// Verilog generated from the al system
`timescale 1ns/10ps
module sine(v,sv);
  input [12:0] v;
  output [15:0] sv;
  reg [15:0] _o_sv;
  assign sv=_o_sv;
  integer _ix_;
  always @(*) begin
    case(v)
      1'b0:
        _o_sv = 1'b0;
      1'b1:
        _o_sv = 3'b110;
      2'b10:
        _o_sv = 4'b1100;
      2'b11:
        _o_sv = 5'b10010;
      3'b100:
        _o_sv = 5'b11001;
      3'b101:
        _o_sv = 5'b11111;
      3'b110:
        _o_sv = 6'b100101;
      3'b111:
        _o_sv = 6'b101011;
      4'b1000:
        _o_sv = 6'b110010;
      4'b1001:
        _o_sv = 6'b111000;
      4'b1010:
        _o_sv = 6'b111110;
      4'b1011:
        _o_sv = 7'b1000101;
      4'b1100:
        _o_sv = 7'b1001011;
      4'b1101:
        _o_sv = 7'b1010001;
      4'b1110:
        _o_sv = 7'b1010111;
      4'b1111:
        _o_sv = 7'b1011110;
      5'b10000:
        _o_sv = 7'b1100100;
      5'b10001:
        _o_sv = 7'b1101010;
      5'b10010:
        _o_sv = 7'b1110001;
      5'b10011:
        _o_sv = 7'b1110111;
      5'b10100:
        _o_sv = 7'b1111101;
      5'b10101:
        _o_sv = 8'b10000011;
      5'b10110:
        _o_sv = 8'b10001010;
      5'b10111:
        _o_sv = 8'b10010000;
      5'b11000:
        _o_sv = 8'b10010110;
      5'b11001:
        _o_sv = 8'b10011101;
      5'b11010:
        _o_sv = 8'b10100011;
      5'b11011:
        _o_sv = 8'b10101001;
      5'b11100:
        _o_sv = 8'b10101111;
      5'b11101:
        _o_sv = 8'b10110110;
      5'b11110:
        _o_sv = 8'b10111100;
      5'b11111:
        _o_sv = 8'b11000010;
      6'b100000:
        _o_sv = 8'b11001001;
      6'b100001:
        _o_sv = 8'b11001111;
      6'b100010:
        _o_sv = 8'b11010101;
      6'b100011:
        _o_sv = 8'b11011011;
      6'b100100:
        _o_sv = 8'b11100010;
      6'b100101:
        _o_sv = 8'b11101000;
      6'b100110:
        _o_sv = 8'b11101110;
      6'b100111:
        _o_sv = 8'b11110101;
      6'b101000:
        _o_sv = 8'b11111011;
      6'b101001:
        _o_sv = 9'b100000001;
      6'b101010:
        _o_sv = 9'b100000111;
      6'b101011:
        _o_sv = 9'b100001110;
      6'b101100:
        _o_sv = 9'b100010100;
      6'b101101:
        _o_sv = 9'b100011010;
      6'b101110:
        _o_sv = 9'b100100001;
      6'b101111:
        _o_sv = 9'b100100111;
      6'b110000:
        _o_sv = 9'b100101101;
      6'b110001:
        _o_sv = 9'b100110011;
      6'b110010:
        _o_sv = 9'b100111010;
      6'b110011:
        _o_sv = 9'b101000000;
      6'b110100:
        _o_sv = 9'b101000110;
      6'b110101:
        _o_sv = 9'b101001101;
      6'b110110:
        _o_sv = 9'b101010011;
      6'b110111:
        _o_sv = 9'b101011001;
      6'b111000:
        _o_sv = 9'b101011111;
      6'b111001:
        _o_sv = 9'b101100110;
      6'b111010:
        _o_sv = 9'b101101100;
      6'b111011:
        _o_sv = 9'b101110010;
      6'b111100:
        _o_sv = 9'b101111000;
      6'b111101:
        _o_sv = 9'b101111111;
      6'b111110:
        _o_sv = 9'b110000101;
      6'b111111:
        _o_sv = 9'b110001011;
      7'b1000000:
        _o_sv = 9'b110010010;
      7'b1000001:
        _o_sv = 9'b110011000;
      7'b1000010:
        _o_sv = 9'b110011110;
      7'b1000011:
        _o_sv = 9'b110100100;
      7'b1000100:
        _o_sv = 9'b110101011;
      7'b1000101:
        _o_sv = 9'b110110001;
      7'b1000110:
        _o_sv = 9'b110110111;
      7'b1000111:
        _o_sv = 9'b110111110;
      7'b1001000:
        _o_sv = 9'b111000100;
      7'b1001001:
        _o_sv = 9'b111001010;
      7'b1001010:
        _o_sv = 9'b111010000;
      7'b1001011:
        _o_sv = 9'b111010111;
      7'b1001100:
        _o_sv = 9'b111011101;
      7'b1001101:
        _o_sv = 9'b111100011;
      7'b1001110:
        _o_sv = 9'b111101010;
      7'b1001111:
        _o_sv = 9'b111110000;
      7'b1010000:
        _o_sv = 9'b111110110;
      7'b1010001:
        _o_sv = 9'b111111100;
      7'b1010010:
        _o_sv = 10'b1000000011;
      7'b1010011:
        _o_sv = 10'b1000001001;
      7'b1010100:
        _o_sv = 10'b1000001111;
      7'b1010101:
        _o_sv = 10'b1000010110;
      7'b1010110:
        _o_sv = 10'b1000011100;
      7'b1010111:
        _o_sv = 10'b1000100010;
      7'b1011000:
        _o_sv = 10'b1000101000;
      7'b1011001:
        _o_sv = 10'b1000101111;
      7'b1011010:
        _o_sv = 10'b1000110101;
      7'b1011011:
        _o_sv = 10'b1000111011;
      7'b1011100:
        _o_sv = 10'b1001000010;
      7'b1011101:
        _o_sv = 10'b1001001000;
      7'b1011110:
        _o_sv = 10'b1001001110;
      7'b1011111:
        _o_sv = 10'b1001010100;
      7'b1100000:
        _o_sv = 10'b1001011011;
      7'b1100001:
        _o_sv = 10'b1001100001;
      7'b1100010:
        _o_sv = 10'b1001100111;
      7'b1100011:
        _o_sv = 10'b1001101101;
      7'b1100100:
        _o_sv = 10'b1001110100;
      7'b1100101:
        _o_sv = 10'b1001111010;
      7'b1100110:
        _o_sv = 10'b1010000000;
      7'b1100111:
        _o_sv = 10'b1010000111;
      7'b1101000:
        _o_sv = 10'b1010001101;
      7'b1101001:
        _o_sv = 10'b1010010011;
      7'b1101010:
        _o_sv = 10'b1010011001;
      7'b1101011:
        _o_sv = 10'b1010100000;
      7'b1101100:
        _o_sv = 10'b1010100110;
      7'b1101101:
        _o_sv = 10'b1010101100;
      7'b1101110:
        _o_sv = 10'b1010110011;
      7'b1101111:
        _o_sv = 10'b1010111001;
      7'b1110000:
        _o_sv = 10'b1010111111;
      7'b1110001:
        _o_sv = 10'b1011000101;
      7'b1110010:
        _o_sv = 10'b1011001100;
      7'b1110011:
        _o_sv = 10'b1011010010;
      7'b1110100:
        _o_sv = 10'b1011011000;
      7'b1110101:
        _o_sv = 10'b1011011111;
      7'b1110110:
        _o_sv = 10'b1011100101;
      7'b1110111:
        _o_sv = 10'b1011101011;
      7'b1111000:
        _o_sv = 10'b1011110001;
      7'b1111001:
        _o_sv = 10'b1011111000;
      7'b1111010:
        _o_sv = 10'b1011111110;
      7'b1111011:
        _o_sv = 10'b1100000100;
      7'b1111100:
        _o_sv = 10'b1100001011;
      7'b1111101:
        _o_sv = 10'b1100010001;
      7'b1111110:
        _o_sv = 10'b1100010111;
      7'b1111111:
        _o_sv = 10'b1100011101;
      8'b10000000:
        _o_sv = 10'b1100100100;
      8'b10000001:
        _o_sv = 10'b1100101010;
      8'b10000010:
        _o_sv = 10'b1100110000;
      8'b10000011:
        _o_sv = 10'b1100110111;
      8'b10000100:
        _o_sv = 10'b1100111101;
      8'b10000101:
        _o_sv = 10'b1101000011;
      8'b10000110:
        _o_sv = 10'b1101001001;
      8'b10000111:
        _o_sv = 10'b1101010000;
      8'b10001000:
        _o_sv = 10'b1101010110;
      8'b10001001:
        _o_sv = 10'b1101011100;
      8'b10001010:
        _o_sv = 10'b1101100010;
      8'b10001011:
        _o_sv = 10'b1101101001;
      8'b10001100:
        _o_sv = 10'b1101101111;
      8'b10001101:
        _o_sv = 10'b1101110101;
      8'b10001110:
        _o_sv = 10'b1101111100;
      8'b10001111:
        _o_sv = 10'b1110000010;
      8'b10010000:
        _o_sv = 10'b1110001000;
      8'b10010001:
        _o_sv = 10'b1110001110;
      8'b10010010:
        _o_sv = 10'b1110010101;
      8'b10010011:
        _o_sv = 10'b1110011011;
      8'b10010100:
        _o_sv = 10'b1110100001;
      8'b10010101:
        _o_sv = 10'b1110101000;
      8'b10010110:
        _o_sv = 10'b1110101110;
      8'b10010111:
        _o_sv = 10'b1110110100;
      8'b10011000:
        _o_sv = 10'b1110111010;
      8'b10011001:
        _o_sv = 10'b1111000001;
      8'b10011010:
        _o_sv = 10'b1111000111;
      8'b10011011:
        _o_sv = 10'b1111001101;
      8'b10011100:
        _o_sv = 10'b1111010100;
      8'b10011101:
        _o_sv = 10'b1111011010;
      8'b10011110:
        _o_sv = 10'b1111100000;
      8'b10011111:
        _o_sv = 10'b1111100110;
      8'b10100000:
        _o_sv = 10'b1111101101;
      8'b10100001:
        _o_sv = 10'b1111110011;
      8'b10100010:
        _o_sv = 10'b1111111001;
      8'b10100011:
        _o_sv = 10'b1111111111;
      8'b10100100:
        _o_sv = 11'b10000000110;
      8'b10100101:
        _o_sv = 11'b10000001100;
      8'b10100110:
        _o_sv = 11'b10000010010;
      8'b10100111:
        _o_sv = 11'b10000011001;
      8'b10101000:
        _o_sv = 11'b10000011111;
      8'b10101001:
        _o_sv = 11'b10000100101;
      8'b10101010:
        _o_sv = 11'b10000101011;
      8'b10101011:
        _o_sv = 11'b10000110010;
      8'b10101100:
        _o_sv = 11'b10000111000;
      8'b10101101:
        _o_sv = 11'b10000111110;
      8'b10101110:
        _o_sv = 11'b10001000101;
      8'b10101111:
        _o_sv = 11'b10001001011;
      8'b10110000:
        _o_sv = 11'b10001010001;
      8'b10110001:
        _o_sv = 11'b10001010111;
      8'b10110010:
        _o_sv = 11'b10001011110;
      8'b10110011:
        _o_sv = 11'b10001100100;
      8'b10110100:
        _o_sv = 11'b10001101010;
      8'b10110101:
        _o_sv = 11'b10001110001;
      8'b10110110:
        _o_sv = 11'b10001110111;
      8'b10110111:
        _o_sv = 11'b10001111101;
      8'b10111000:
        _o_sv = 11'b10010000011;
      8'b10111001:
        _o_sv = 11'b10010001010;
      8'b10111010:
        _o_sv = 11'b10010010000;
      8'b10111011:
        _o_sv = 11'b10010010110;
      8'b10111100:
        _o_sv = 11'b10010011100;
      8'b10111101:
        _o_sv = 11'b10010100011;
      8'b10111110:
        _o_sv = 11'b10010101001;
      8'b10111111:
        _o_sv = 11'b10010101111;
      8'b11000000:
        _o_sv = 11'b10010110110;
      8'b11000001:
        _o_sv = 11'b10010111100;
      8'b11000010:
        _o_sv = 11'b10011000010;
      8'b11000011:
        _o_sv = 11'b10011001000;
      8'b11000100:
        _o_sv = 11'b10011001111;
      8'b11000101:
        _o_sv = 11'b10011010101;
      8'b11000110:
        _o_sv = 11'b10011011011;
      8'b11000111:
        _o_sv = 11'b10011100010;
      8'b11001000:
        _o_sv = 11'b10011101000;
      8'b11001001:
        _o_sv = 11'b10011101110;
      8'b11001010:
        _o_sv = 11'b10011110100;
      8'b11001011:
        _o_sv = 11'b10011111011;
      8'b11001100:
        _o_sv = 11'b10100000001;
      8'b11001101:
        _o_sv = 11'b10100000111;
      8'b11001110:
        _o_sv = 11'b10100001101;
      8'b11001111:
        _o_sv = 11'b10100010100;
      8'b11010000:
        _o_sv = 11'b10100011010;
      8'b11010001:
        _o_sv = 11'b10100100000;
      8'b11010010:
        _o_sv = 11'b10100100111;
      8'b11010011:
        _o_sv = 11'b10100101101;
      8'b11010100:
        _o_sv = 11'b10100110011;
      8'b11010101:
        _o_sv = 11'b10100111001;
      8'b11010110:
        _o_sv = 11'b10101000000;
      8'b11010111:
        _o_sv = 11'b10101000110;
      8'b11011000:
        _o_sv = 11'b10101001100;
      8'b11011001:
        _o_sv = 11'b10101010011;
      8'b11011010:
        _o_sv = 11'b10101011001;
      8'b11011011:
        _o_sv = 11'b10101011111;
      8'b11011100:
        _o_sv = 11'b10101100101;
      8'b11011101:
        _o_sv = 11'b10101101100;
      8'b11011110:
        _o_sv = 11'b10101110010;
      8'b11011111:
        _o_sv = 11'b10101111000;
      8'b11100000:
        _o_sv = 11'b10101111111;
      8'b11100001:
        _o_sv = 11'b10110000101;
      8'b11100010:
        _o_sv = 11'b10110001011;
      8'b11100011:
        _o_sv = 11'b10110010001;
      8'b11100100:
        _o_sv = 11'b10110011000;
      8'b11100101:
        _o_sv = 11'b10110011110;
      8'b11100110:
        _o_sv = 11'b10110100100;
      8'b11100111:
        _o_sv = 11'b10110101010;
      8'b11101000:
        _o_sv = 11'b10110110001;
      8'b11101001:
        _o_sv = 11'b10110110111;
      8'b11101010:
        _o_sv = 11'b10110111101;
      8'b11101011:
        _o_sv = 11'b10111000100;
      8'b11101100:
        _o_sv = 11'b10111001010;
      8'b11101101:
        _o_sv = 11'b10111010000;
      8'b11101110:
        _o_sv = 11'b10111010110;
      8'b11101111:
        _o_sv = 11'b10111011101;
      8'b11110000:
        _o_sv = 11'b10111100011;
      8'b11110001:
        _o_sv = 11'b10111101001;
      8'b11110010:
        _o_sv = 11'b10111101111;
      8'b11110011:
        _o_sv = 11'b10111110110;
      8'b11110100:
        _o_sv = 11'b10111111100;
      8'b11110101:
        _o_sv = 11'b11000000010;
      8'b11110110:
        _o_sv = 11'b11000001001;
      8'b11110111:
        _o_sv = 11'b11000001111;
      8'b11111000:
        _o_sv = 11'b11000010101;
      8'b11111001:
        _o_sv = 11'b11000011011;
      8'b11111010:
        _o_sv = 11'b11000100010;
      8'b11111011:
        _o_sv = 11'b11000101000;
      8'b11111100:
        _o_sv = 11'b11000101110;
      8'b11111101:
        _o_sv = 11'b11000110101;
      8'b11111110:
        _o_sv = 11'b11000111011;
      8'b11111111:
        _o_sv = 11'b11001000001;
      9'b100000000:
        _o_sv = 11'b11001000111;
      9'b100000001:
        _o_sv = 11'b11001001110;
      9'b100000010:
        _o_sv = 11'b11001010100;
      9'b100000011:
        _o_sv = 11'b11001011010;
      9'b100000100:
        _o_sv = 11'b11001100000;
      9'b100000101:
        _o_sv = 11'b11001100111;
      9'b100000110:
        _o_sv = 11'b11001101101;
      9'b100000111:
        _o_sv = 11'b11001110011;
      9'b100001000:
        _o_sv = 11'b11001111010;
      9'b100001001:
        _o_sv = 11'b11010000000;
      9'b100001010:
        _o_sv = 11'b11010000110;
      9'b100001011:
        _o_sv = 11'b11010001100;
      9'b100001100:
        _o_sv = 11'b11010010011;
      9'b100001101:
        _o_sv = 11'b11010011001;
      9'b100001110:
        _o_sv = 11'b11010011111;
      9'b100001111:
        _o_sv = 11'b11010100101;
      9'b100010000:
        _o_sv = 11'b11010101100;
      9'b100010001:
        _o_sv = 11'b11010110010;
      9'b100010010:
        _o_sv = 11'b11010111000;
      9'b100010011:
        _o_sv = 11'b11010111111;
      9'b100010100:
        _o_sv = 11'b11011000101;
      9'b100010101:
        _o_sv = 11'b11011001011;
      9'b100010110:
        _o_sv = 11'b11011010001;
      9'b100010111:
        _o_sv = 11'b11011011000;
      9'b100011000:
        _o_sv = 11'b11011011110;
      9'b100011001:
        _o_sv = 11'b11011100100;
      9'b100011010:
        _o_sv = 11'b11011101010;
      9'b100011011:
        _o_sv = 11'b11011110001;
      9'b100011100:
        _o_sv = 11'b11011110111;
      9'b100011101:
        _o_sv = 11'b11011111101;
      9'b100011110:
        _o_sv = 11'b11100000100;
      9'b100011111:
        _o_sv = 11'b11100001010;
      9'b100100000:
        _o_sv = 11'b11100010000;
      9'b100100001:
        _o_sv = 11'b11100010110;
      9'b100100010:
        _o_sv = 11'b11100011101;
      9'b100100011:
        _o_sv = 11'b11100100011;
      9'b100100100:
        _o_sv = 11'b11100101001;
      9'b100100101:
        _o_sv = 11'b11100110000;
      9'b100100110:
        _o_sv = 11'b11100110110;
      9'b100100111:
        _o_sv = 11'b11100111100;
      9'b100101000:
        _o_sv = 11'b11101000010;
      9'b100101001:
        _o_sv = 11'b11101001001;
      9'b100101010:
        _o_sv = 11'b11101001111;
      9'b100101011:
        _o_sv = 11'b11101010101;
      9'b100101100:
        _o_sv = 11'b11101011011;
      9'b100101101:
        _o_sv = 11'b11101100010;
      9'b100101110:
        _o_sv = 11'b11101101000;
      9'b100101111:
        _o_sv = 11'b11101101110;
      9'b100110000:
        _o_sv = 11'b11101110101;
      9'b100110001:
        _o_sv = 11'b11101111011;
      9'b100110010:
        _o_sv = 11'b11110000001;
      9'b100110011:
        _o_sv = 11'b11110000111;
      9'b100110100:
        _o_sv = 11'b11110001110;
      9'b100110101:
        _o_sv = 11'b11110010100;
      9'b100110110:
        _o_sv = 11'b11110011010;
      9'b100110111:
        _o_sv = 11'b11110100000;
      9'b100111000:
        _o_sv = 11'b11110100111;
      9'b100111001:
        _o_sv = 11'b11110101101;
      9'b100111010:
        _o_sv = 11'b11110110011;
      9'b100111011:
        _o_sv = 11'b11110111010;
      9'b100111100:
        _o_sv = 11'b11111000000;
      9'b100111101:
        _o_sv = 11'b11111000110;
      9'b100111110:
        _o_sv = 11'b11111001100;
      9'b100111111:
        _o_sv = 11'b11111010011;
      9'b101000000:
        _o_sv = 11'b11111011001;
      9'b101000001:
        _o_sv = 11'b11111011111;
      9'b101000010:
        _o_sv = 11'b11111100101;
      9'b101000011:
        _o_sv = 11'b11111101100;
      9'b101000100:
        _o_sv = 11'b11111110010;
      9'b101000101:
        _o_sv = 11'b11111111000;
      9'b101000110:
        _o_sv = 11'b11111111110;
      9'b101000111:
        _o_sv = 12'b100000000101;
      9'b101001000:
        _o_sv = 12'b100000001011;
      9'b101001001:
        _o_sv = 12'b100000010001;
      9'b101001010:
        _o_sv = 12'b100000011000;
      9'b101001011:
        _o_sv = 12'b100000011110;
      9'b101001100:
        _o_sv = 12'b100000100100;
      9'b101001101:
        _o_sv = 12'b100000101010;
      9'b101001110:
        _o_sv = 12'b100000110001;
      9'b101001111:
        _o_sv = 12'b100000110111;
      9'b101010000:
        _o_sv = 12'b100000111101;
      9'b101010001:
        _o_sv = 12'b100001000011;
      9'b101010010:
        _o_sv = 12'b100001001010;
      9'b101010011:
        _o_sv = 12'b100001010000;
      9'b101010100:
        _o_sv = 12'b100001010110;
      9'b101010101:
        _o_sv = 12'b100001011101;
      9'b101010110:
        _o_sv = 12'b100001100011;
      9'b101010111:
        _o_sv = 12'b100001101001;
      9'b101011000:
        _o_sv = 12'b100001101111;
      9'b101011001:
        _o_sv = 12'b100001110110;
      9'b101011010:
        _o_sv = 12'b100001111100;
      9'b101011011:
        _o_sv = 12'b100010000010;
      9'b101011100:
        _o_sv = 12'b100010001000;
      9'b101011101:
        _o_sv = 12'b100010001111;
      9'b101011110:
        _o_sv = 12'b100010010101;
      9'b101011111:
        _o_sv = 12'b100010011011;
      9'b101100000:
        _o_sv = 12'b100010100010;
      9'b101100001:
        _o_sv = 12'b100010101000;
      9'b101100010:
        _o_sv = 12'b100010101110;
      9'b101100011:
        _o_sv = 12'b100010110100;
      9'b101100100:
        _o_sv = 12'b100010111011;
      9'b101100101:
        _o_sv = 12'b100011000001;
      9'b101100110:
        _o_sv = 12'b100011000111;
      9'b101100111:
        _o_sv = 12'b100011001101;
      9'b101101000:
        _o_sv = 12'b100011010100;
      9'b101101001:
        _o_sv = 12'b100011011010;
      9'b101101010:
        _o_sv = 12'b100011100000;
      9'b101101011:
        _o_sv = 12'b100011100110;
      9'b101101100:
        _o_sv = 12'b100011101101;
      9'b101101101:
        _o_sv = 12'b100011110011;
      9'b101101110:
        _o_sv = 12'b100011111001;
      9'b101101111:
        _o_sv = 12'b100100000000;
      9'b101110000:
        _o_sv = 12'b100100000110;
      9'b101110001:
        _o_sv = 12'b100100001100;
      9'b101110010:
        _o_sv = 12'b100100010010;
      9'b101110011:
        _o_sv = 12'b100100011001;
      9'b101110100:
        _o_sv = 12'b100100011111;
      9'b101110101:
        _o_sv = 12'b100100100101;
      9'b101110110:
        _o_sv = 12'b100100101011;
      9'b101110111:
        _o_sv = 12'b100100110010;
      9'b101111000:
        _o_sv = 12'b100100111000;
      9'b101111001:
        _o_sv = 12'b100100111110;
      9'b101111010:
        _o_sv = 12'b100101000100;
      9'b101111011:
        _o_sv = 12'b100101001011;
      9'b101111100:
        _o_sv = 12'b100101010001;
      9'b101111101:
        _o_sv = 12'b100101010111;
      9'b101111110:
        _o_sv = 12'b100101011110;
      9'b101111111:
        _o_sv = 12'b100101100100;
      9'b110000000:
        _o_sv = 12'b100101101010;
      9'b110000001:
        _o_sv = 12'b100101110000;
      9'b110000010:
        _o_sv = 12'b100101110111;
      9'b110000011:
        _o_sv = 12'b100101111101;
      9'b110000100:
        _o_sv = 12'b100110000011;
      9'b110000101:
        _o_sv = 12'b100110001001;
      9'b110000110:
        _o_sv = 12'b100110010000;
      9'b110000111:
        _o_sv = 12'b100110010110;
      9'b110001000:
        _o_sv = 12'b100110011100;
      9'b110001001:
        _o_sv = 12'b100110100010;
      9'b110001010:
        _o_sv = 12'b100110101001;
      9'b110001011:
        _o_sv = 12'b100110101111;
      9'b110001100:
        _o_sv = 12'b100110110101;
      9'b110001101:
        _o_sv = 12'b100110111100;
      9'b110001110:
        _o_sv = 12'b100111000010;
      9'b110001111:
        _o_sv = 12'b100111001000;
      9'b110010000:
        _o_sv = 12'b100111001110;
      9'b110010001:
        _o_sv = 12'b100111010101;
      9'b110010010:
        _o_sv = 12'b100111011011;
      9'b110010011:
        _o_sv = 12'b100111100001;
      9'b110010100:
        _o_sv = 12'b100111100111;
      9'b110010101:
        _o_sv = 12'b100111101110;
      9'b110010110:
        _o_sv = 12'b100111110100;
      9'b110010111:
        _o_sv = 12'b100111111010;
      9'b110011000:
        _o_sv = 12'b101000000000;
      9'b110011001:
        _o_sv = 12'b101000000111;
      9'b110011010:
        _o_sv = 12'b101000001101;
      9'b110011011:
        _o_sv = 12'b101000010011;
      9'b110011100:
        _o_sv = 12'b101000011001;
      9'b110011101:
        _o_sv = 12'b101000100000;
      9'b110011110:
        _o_sv = 12'b101000100110;
      9'b110011111:
        _o_sv = 12'b101000101100;
      9'b110100000:
        _o_sv = 12'b101000110011;
      9'b110100001:
        _o_sv = 12'b101000111001;
      9'b110100010:
        _o_sv = 12'b101000111111;
      9'b110100011:
        _o_sv = 12'b101001000101;
      9'b110100100:
        _o_sv = 12'b101001001100;
      9'b110100101:
        _o_sv = 12'b101001010010;
      9'b110100110:
        _o_sv = 12'b101001011000;
      9'b110100111:
        _o_sv = 12'b101001011110;
      9'b110101000:
        _o_sv = 12'b101001100101;
      9'b110101001:
        _o_sv = 12'b101001101011;
      9'b110101010:
        _o_sv = 12'b101001110001;
      9'b110101011:
        _o_sv = 12'b101001110111;
      9'b110101100:
        _o_sv = 12'b101001111110;
      9'b110101101:
        _o_sv = 12'b101010000100;
      9'b110101110:
        _o_sv = 12'b101010001010;
      9'b110101111:
        _o_sv = 12'b101010010000;
      9'b110110000:
        _o_sv = 12'b101010010111;
      9'b110110001:
        _o_sv = 12'b101010011101;
      9'b110110010:
        _o_sv = 12'b101010100011;
      9'b110110011:
        _o_sv = 12'b101010101010;
      9'b110110100:
        _o_sv = 12'b101010110000;
      9'b110110101:
        _o_sv = 12'b101010110110;
      9'b110110110:
        _o_sv = 12'b101010111100;
      9'b110110111:
        _o_sv = 12'b101011000011;
      9'b110111000:
        _o_sv = 12'b101011001001;
      9'b110111001:
        _o_sv = 12'b101011001111;
      9'b110111010:
        _o_sv = 12'b101011010101;
      9'b110111011:
        _o_sv = 12'b101011011100;
      9'b110111100:
        _o_sv = 12'b101011100010;
      9'b110111101:
        _o_sv = 12'b101011101000;
      9'b110111110:
        _o_sv = 12'b101011101110;
      9'b110111111:
        _o_sv = 12'b101011110101;
      9'b111000000:
        _o_sv = 12'b101011111011;
      9'b111000001:
        _o_sv = 12'b101100000001;
      9'b111000010:
        _o_sv = 12'b101100000111;
      9'b111000011:
        _o_sv = 12'b101100001110;
      9'b111000100:
        _o_sv = 12'b101100010100;
      9'b111000101:
        _o_sv = 12'b101100011010;
      9'b111000110:
        _o_sv = 12'b101100100000;
      9'b111000111:
        _o_sv = 12'b101100100111;
      9'b111001000:
        _o_sv = 12'b101100101101;
      9'b111001001:
        _o_sv = 12'b101100110011;
      9'b111001010:
        _o_sv = 12'b101100111010;
      9'b111001011:
        _o_sv = 12'b101101000000;
      9'b111001100:
        _o_sv = 12'b101101000110;
      9'b111001101:
        _o_sv = 12'b101101001100;
      9'b111001110:
        _o_sv = 12'b101101010011;
      9'b111001111:
        _o_sv = 12'b101101011001;
      9'b111010000:
        _o_sv = 12'b101101011111;
      9'b111010001:
        _o_sv = 12'b101101100101;
      9'b111010010:
        _o_sv = 12'b101101101100;
      9'b111010011:
        _o_sv = 12'b101101110010;
      9'b111010100:
        _o_sv = 12'b101101111000;
      9'b111010101:
        _o_sv = 12'b101101111110;
      9'b111010110:
        _o_sv = 12'b101110000101;
      9'b111010111:
        _o_sv = 12'b101110001011;
      9'b111011000:
        _o_sv = 12'b101110010001;
      9'b111011001:
        _o_sv = 12'b101110010111;
      9'b111011010:
        _o_sv = 12'b101110011110;
      9'b111011011:
        _o_sv = 12'b101110100100;
      9'b111011100:
        _o_sv = 12'b101110101010;
      9'b111011101:
        _o_sv = 12'b101110110000;
      9'b111011110:
        _o_sv = 12'b101110110111;
      9'b111011111:
        _o_sv = 12'b101110111101;
      9'b111100000:
        _o_sv = 12'b101111000011;
      9'b111100001:
        _o_sv = 12'b101111001001;
      9'b111100010:
        _o_sv = 12'b101111010000;
      9'b111100011:
        _o_sv = 12'b101111010110;
      9'b111100100:
        _o_sv = 12'b101111011100;
      9'b111100101:
        _o_sv = 12'b101111100010;
      9'b111100110:
        _o_sv = 12'b101111101001;
      9'b111100111:
        _o_sv = 12'b101111101111;
      9'b111101000:
        _o_sv = 12'b101111110101;
      9'b111101001:
        _o_sv = 12'b101111111011;
      9'b111101010:
        _o_sv = 12'b110000000010;
      9'b111101011:
        _o_sv = 12'b110000001000;
      9'b111101100:
        _o_sv = 12'b110000001110;
      9'b111101101:
        _o_sv = 12'b110000010100;
      9'b111101110:
        _o_sv = 12'b110000011011;
      9'b111101111:
        _o_sv = 12'b110000100001;
      9'b111110000:
        _o_sv = 12'b110000100111;
      9'b111110001:
        _o_sv = 12'b110000101110;
      9'b111110010:
        _o_sv = 12'b110000110100;
      9'b111110011:
        _o_sv = 12'b110000111010;
      9'b111110100:
        _o_sv = 12'b110001000000;
      9'b111110101:
        _o_sv = 12'b110001000111;
      9'b111110110:
        _o_sv = 12'b110001001101;
      9'b111110111:
        _o_sv = 12'b110001010011;
      9'b111111000:
        _o_sv = 12'b110001011001;
      9'b111111001:
        _o_sv = 12'b110001100000;
      9'b111111010:
        _o_sv = 12'b110001100110;
      9'b111111011:
        _o_sv = 12'b110001101100;
      9'b111111100:
        _o_sv = 12'b110001110010;
      9'b111111101:
        _o_sv = 12'b110001111001;
      9'b111111110:
        _o_sv = 12'b110001111111;
      9'b111111111:
        _o_sv = 12'b110010000101;
      10'b1000000000:
        _o_sv = 12'b110010001011;
      10'b1000000001:
        _o_sv = 12'b110010010010;
      10'b1000000010:
        _o_sv = 12'b110010011000;
      10'b1000000011:
        _o_sv = 12'b110010011110;
      10'b1000000100:
        _o_sv = 12'b110010100100;
      10'b1000000101:
        _o_sv = 12'b110010101011;
      10'b1000000110:
        _o_sv = 12'b110010110001;
      10'b1000000111:
        _o_sv = 12'b110010110111;
      10'b1000001000:
        _o_sv = 12'b110010111101;
      10'b1000001001:
        _o_sv = 12'b110011000100;
      10'b1000001010:
        _o_sv = 12'b110011001010;
      10'b1000001011:
        _o_sv = 12'b110011010000;
      10'b1000001100:
        _o_sv = 12'b110011010110;
      10'b1000001101:
        _o_sv = 12'b110011011101;
      10'b1000001110:
        _o_sv = 12'b110011100011;
      10'b1000001111:
        _o_sv = 12'b110011101001;
      10'b1000010000:
        _o_sv = 12'b110011101111;
      10'b1000010001:
        _o_sv = 12'b110011110110;
      10'b1000010010:
        _o_sv = 12'b110011111100;
      10'b1000010011:
        _o_sv = 12'b110100000010;
      10'b1000010100:
        _o_sv = 12'b110100001000;
      10'b1000010101:
        _o_sv = 12'b110100001111;
      10'b1000010110:
        _o_sv = 12'b110100010101;
      10'b1000010111:
        _o_sv = 12'b110100011011;
      10'b1000011000:
        _o_sv = 12'b110100100001;
      10'b1000011001:
        _o_sv = 12'b110100101000;
      10'b1000011010:
        _o_sv = 12'b110100101110;
      10'b1000011011:
        _o_sv = 12'b110100110100;
      10'b1000011100:
        _o_sv = 12'b110100111010;
      10'b1000011101:
        _o_sv = 12'b110101000001;
      10'b1000011110:
        _o_sv = 12'b110101000111;
      10'b1000011111:
        _o_sv = 12'b110101001101;
      10'b1000100000:
        _o_sv = 12'b110101010011;
      10'b1000100001:
        _o_sv = 12'b110101011010;
      10'b1000100010:
        _o_sv = 12'b110101100000;
      10'b1000100011:
        _o_sv = 12'b110101100110;
      10'b1000100100:
        _o_sv = 12'b110101101100;
      10'b1000100101:
        _o_sv = 12'b110101110011;
      10'b1000100110:
        _o_sv = 12'b110101111001;
      10'b1000100111:
        _o_sv = 12'b110101111111;
      10'b1000101000:
        _o_sv = 12'b110110000101;
      10'b1000101001:
        _o_sv = 12'b110110001100;
      10'b1000101010:
        _o_sv = 12'b110110010010;
      10'b1000101011:
        _o_sv = 12'b110110011000;
      10'b1000101100:
        _o_sv = 12'b110110011110;
      10'b1000101101:
        _o_sv = 12'b110110100101;
      10'b1000101110:
        _o_sv = 12'b110110101011;
      10'b1000101111:
        _o_sv = 12'b110110110001;
      10'b1000110000:
        _o_sv = 12'b110110110111;
      10'b1000110001:
        _o_sv = 12'b110110111110;
      10'b1000110010:
        _o_sv = 12'b110111000100;
      10'b1000110011:
        _o_sv = 12'b110111001010;
      10'b1000110100:
        _o_sv = 12'b110111010000;
      10'b1000110101:
        _o_sv = 12'b110111010111;
      10'b1000110110:
        _o_sv = 12'b110111011101;
      10'b1000110111:
        _o_sv = 12'b110111100011;
      10'b1000111000:
        _o_sv = 12'b110111101001;
      10'b1000111001:
        _o_sv = 12'b110111110000;
      10'b1000111010:
        _o_sv = 12'b110111110110;
      10'b1000111011:
        _o_sv = 12'b110111111100;
      10'b1000111100:
        _o_sv = 12'b111000000010;
      10'b1000111101:
        _o_sv = 12'b111000001001;
      10'b1000111110:
        _o_sv = 12'b111000001111;
      10'b1000111111:
        _o_sv = 12'b111000010101;
      10'b1001000000:
        _o_sv = 12'b111000011011;
      10'b1001000001:
        _o_sv = 12'b111000100010;
      10'b1001000010:
        _o_sv = 12'b111000101000;
      10'b1001000011:
        _o_sv = 12'b111000101110;
      10'b1001000100:
        _o_sv = 12'b111000110100;
      10'b1001000101:
        _o_sv = 12'b111000111010;
      10'b1001000110:
        _o_sv = 12'b111001000001;
      10'b1001000111:
        _o_sv = 12'b111001000111;
      10'b1001001000:
        _o_sv = 12'b111001001101;
      10'b1001001001:
        _o_sv = 12'b111001010011;
      10'b1001001010:
        _o_sv = 12'b111001011010;
      10'b1001001011:
        _o_sv = 12'b111001100000;
      10'b1001001100:
        _o_sv = 12'b111001100110;
      10'b1001001101:
        _o_sv = 12'b111001101100;
      10'b1001001110:
        _o_sv = 12'b111001110011;
      10'b1001001111:
        _o_sv = 12'b111001111001;
      10'b1001010000:
        _o_sv = 12'b111001111111;
      10'b1001010001:
        _o_sv = 12'b111010000101;
      10'b1001010010:
        _o_sv = 12'b111010001100;
      10'b1001010011:
        _o_sv = 12'b111010010010;
      10'b1001010100:
        _o_sv = 12'b111010011000;
      10'b1001010101:
        _o_sv = 12'b111010011110;
      10'b1001010110:
        _o_sv = 12'b111010100101;
      10'b1001010111:
        _o_sv = 12'b111010101011;
      10'b1001011000:
        _o_sv = 12'b111010110001;
      10'b1001011001:
        _o_sv = 12'b111010110111;
      10'b1001011010:
        _o_sv = 12'b111010111110;
      10'b1001011011:
        _o_sv = 12'b111011000100;
      10'b1001011100:
        _o_sv = 12'b111011001010;
      10'b1001011101:
        _o_sv = 12'b111011010000;
      10'b1001011110:
        _o_sv = 12'b111011010111;
      10'b1001011111:
        _o_sv = 12'b111011011101;
      10'b1001100000:
        _o_sv = 12'b111011100011;
      10'b1001100001:
        _o_sv = 12'b111011101001;
      10'b1001100010:
        _o_sv = 12'b111011110000;
      10'b1001100011:
        _o_sv = 12'b111011110110;
      10'b1001100100:
        _o_sv = 12'b111011111100;
      10'b1001100101:
        _o_sv = 12'b111100000010;
      10'b1001100110:
        _o_sv = 12'b111100001000;
      10'b1001100111:
        _o_sv = 12'b111100001111;
      10'b1001101000:
        _o_sv = 12'b111100010101;
      10'b1001101001:
        _o_sv = 12'b111100011011;
      10'b1001101010:
        _o_sv = 12'b111100100001;
      10'b1001101011:
        _o_sv = 12'b111100101000;
      10'b1001101100:
        _o_sv = 12'b111100101110;
      10'b1001101101:
        _o_sv = 12'b111100110100;
      10'b1001101110:
        _o_sv = 12'b111100111010;
      10'b1001101111:
        _o_sv = 12'b111101000001;
      10'b1001110000:
        _o_sv = 12'b111101000111;
      10'b1001110001:
        _o_sv = 12'b111101001101;
      10'b1001110010:
        _o_sv = 12'b111101010011;
      10'b1001110011:
        _o_sv = 12'b111101011010;
      10'b1001110100:
        _o_sv = 12'b111101100000;
      10'b1001110101:
        _o_sv = 12'b111101100110;
      10'b1001110110:
        _o_sv = 12'b111101101100;
      10'b1001110111:
        _o_sv = 12'b111101110011;
      10'b1001111000:
        _o_sv = 12'b111101111001;
      10'b1001111001:
        _o_sv = 12'b111101111111;
      10'b1001111010:
        _o_sv = 12'b111110000101;
      10'b1001111011:
        _o_sv = 12'b111110001011;
      10'b1001111100:
        _o_sv = 12'b111110010010;
      10'b1001111101:
        _o_sv = 12'b111110011000;
      10'b1001111110:
        _o_sv = 12'b111110011110;
      10'b1001111111:
        _o_sv = 12'b111110100100;
      10'b1010000000:
        _o_sv = 12'b111110101011;
      10'b1010000001:
        _o_sv = 12'b111110110001;
      10'b1010000010:
        _o_sv = 12'b111110110111;
      10'b1010000011:
        _o_sv = 12'b111110111101;
      10'b1010000100:
        _o_sv = 12'b111111000100;
      10'b1010000101:
        _o_sv = 12'b111111001010;
      10'b1010000110:
        _o_sv = 12'b111111010000;
      10'b1010000111:
        _o_sv = 12'b111111010110;
      10'b1010001000:
        _o_sv = 12'b111111011101;
      10'b1010001001:
        _o_sv = 12'b111111100011;
      10'b1010001010:
        _o_sv = 12'b111111101001;
      10'b1010001011:
        _o_sv = 12'b111111101111;
      10'b1010001100:
        _o_sv = 12'b111111110101;
      10'b1010001101:
        _o_sv = 12'b111111111100;
      10'b1010001110:
        _o_sv = 13'b1000000000010;
      10'b1010001111:
        _o_sv = 13'b1000000001000;
      10'b1010010000:
        _o_sv = 13'b1000000001110;
      10'b1010010001:
        _o_sv = 13'b1000000010101;
      10'b1010010010:
        _o_sv = 13'b1000000011011;
      10'b1010010011:
        _o_sv = 13'b1000000100001;
      10'b1010010100:
        _o_sv = 13'b1000000100111;
      10'b1010010101:
        _o_sv = 13'b1000000101110;
      10'b1010010110:
        _o_sv = 13'b1000000110100;
      10'b1010010111:
        _o_sv = 13'b1000000111010;
      10'b1010011000:
        _o_sv = 13'b1000001000000;
      10'b1010011001:
        _o_sv = 13'b1000001000111;
      10'b1010011010:
        _o_sv = 13'b1000001001101;
      10'b1010011011:
        _o_sv = 13'b1000001010011;
      10'b1010011100:
        _o_sv = 13'b1000001011001;
      10'b1010011101:
        _o_sv = 13'b1000001011111;
      10'b1010011110:
        _o_sv = 13'b1000001100110;
      10'b1010011111:
        _o_sv = 13'b1000001101100;
      10'b1010100000:
        _o_sv = 13'b1000001110010;
      10'b1010100001:
        _o_sv = 13'b1000001111000;
      10'b1010100010:
        _o_sv = 13'b1000001111111;
      10'b1010100011:
        _o_sv = 13'b1000010000101;
      10'b1010100100:
        _o_sv = 13'b1000010001011;
      10'b1010100101:
        _o_sv = 13'b1000010010001;
      10'b1010100110:
        _o_sv = 13'b1000010011000;
      10'b1010100111:
        _o_sv = 13'b1000010011110;
      10'b1010101000:
        _o_sv = 13'b1000010100100;
      10'b1010101001:
        _o_sv = 13'b1000010101010;
      10'b1010101010:
        _o_sv = 13'b1000010110000;
      10'b1010101011:
        _o_sv = 13'b1000010110111;
      10'b1010101100:
        _o_sv = 13'b1000010111101;
      10'b1010101101:
        _o_sv = 13'b1000011000011;
      10'b1010101110:
        _o_sv = 13'b1000011001001;
      10'b1010101111:
        _o_sv = 13'b1000011010000;
      10'b1010110000:
        _o_sv = 13'b1000011010110;
      10'b1010110001:
        _o_sv = 13'b1000011011100;
      10'b1010110010:
        _o_sv = 13'b1000011100010;
      10'b1010110011:
        _o_sv = 13'b1000011101000;
      10'b1010110100:
        _o_sv = 13'b1000011101111;
      10'b1010110101:
        _o_sv = 13'b1000011110101;
      10'b1010110110:
        _o_sv = 13'b1000011111011;
      10'b1010110111:
        _o_sv = 13'b1000100000001;
      10'b1010111000:
        _o_sv = 13'b1000100001000;
      10'b1010111001:
        _o_sv = 13'b1000100001110;
      10'b1010111010:
        _o_sv = 13'b1000100010100;
      10'b1010111011:
        _o_sv = 13'b1000100011010;
      10'b1010111100:
        _o_sv = 13'b1000100100001;
      10'b1010111101:
        _o_sv = 13'b1000100100111;
      10'b1010111110:
        _o_sv = 13'b1000100101101;
      10'b1010111111:
        _o_sv = 13'b1000100110011;
      10'b1011000000:
        _o_sv = 13'b1000100111001;
      10'b1011000001:
        _o_sv = 13'b1000101000000;
      10'b1011000010:
        _o_sv = 13'b1000101000110;
      10'b1011000011:
        _o_sv = 13'b1000101001100;
      10'b1011000100:
        _o_sv = 13'b1000101010010;
      10'b1011000101:
        _o_sv = 13'b1000101011001;
      10'b1011000110:
        _o_sv = 13'b1000101011111;
      10'b1011000111:
        _o_sv = 13'b1000101100101;
      10'b1011001000:
        _o_sv = 13'b1000101101011;
      10'b1011001001:
        _o_sv = 13'b1000101110001;
      10'b1011001010:
        _o_sv = 13'b1000101111000;
      10'b1011001011:
        _o_sv = 13'b1000101111110;
      10'b1011001100:
        _o_sv = 13'b1000110000100;
      10'b1011001101:
        _o_sv = 13'b1000110001010;
      10'b1011001110:
        _o_sv = 13'b1000110010001;
      10'b1011001111:
        _o_sv = 13'b1000110010111;
      10'b1011010000:
        _o_sv = 13'b1000110011101;
      10'b1011010001:
        _o_sv = 13'b1000110100011;
      10'b1011010010:
        _o_sv = 13'b1000110101001;
      10'b1011010011:
        _o_sv = 13'b1000110110000;
      10'b1011010100:
        _o_sv = 13'b1000110110110;
      10'b1011010101:
        _o_sv = 13'b1000110111100;
      10'b1011010110:
        _o_sv = 13'b1000111000010;
      10'b1011010111:
        _o_sv = 13'b1000111001001;
      10'b1011011000:
        _o_sv = 13'b1000111001111;
      10'b1011011001:
        _o_sv = 13'b1000111010101;
      10'b1011011010:
        _o_sv = 13'b1000111011011;
      10'b1011011011:
        _o_sv = 13'b1000111100001;
      10'b1011011100:
        _o_sv = 13'b1000111101000;
      10'b1011011101:
        _o_sv = 13'b1000111101110;
      10'b1011011110:
        _o_sv = 13'b1000111110100;
      10'b1011011111:
        _o_sv = 13'b1000111111010;
      10'b1011100000:
        _o_sv = 13'b1001000000001;
      10'b1011100001:
        _o_sv = 13'b1001000000111;
      10'b1011100010:
        _o_sv = 13'b1001000001101;
      10'b1011100011:
        _o_sv = 13'b1001000010011;
      10'b1011100100:
        _o_sv = 13'b1001000011001;
      10'b1011100101:
        _o_sv = 13'b1001000100000;
      10'b1011100110:
        _o_sv = 13'b1001000100110;
      10'b1011100111:
        _o_sv = 13'b1001000101100;
      10'b1011101000:
        _o_sv = 13'b1001000110010;
      10'b1011101001:
        _o_sv = 13'b1001000111001;
      10'b1011101010:
        _o_sv = 13'b1001000111111;
      10'b1011101011:
        _o_sv = 13'b1001001000101;
      10'b1011101100:
        _o_sv = 13'b1001001001011;
      10'b1011101101:
        _o_sv = 13'b1001001010001;
      10'b1011101110:
        _o_sv = 13'b1001001011000;
      10'b1011101111:
        _o_sv = 13'b1001001011110;
      10'b1011110000:
        _o_sv = 13'b1001001100100;
      10'b1011110001:
        _o_sv = 13'b1001001101010;
      10'b1011110010:
        _o_sv = 13'b1001001110001;
      10'b1011110011:
        _o_sv = 13'b1001001110111;
      10'b1011110100:
        _o_sv = 13'b1001001111101;
      10'b1011110101:
        _o_sv = 13'b1001010000011;
      10'b1011110110:
        _o_sv = 13'b1001010001001;
      10'b1011110111:
        _o_sv = 13'b1001010010000;
      10'b1011111000:
        _o_sv = 13'b1001010010110;
      10'b1011111001:
        _o_sv = 13'b1001010011100;
      10'b1011111010:
        _o_sv = 13'b1001010100010;
      10'b1011111011:
        _o_sv = 13'b1001010101000;
      10'b1011111100:
        _o_sv = 13'b1001010101111;
      10'b1011111101:
        _o_sv = 13'b1001010110101;
      10'b1011111110:
        _o_sv = 13'b1001010111011;
      10'b1011111111:
        _o_sv = 13'b1001011000001;
      10'b1100000000:
        _o_sv = 13'b1001011001000;
      10'b1100000001:
        _o_sv = 13'b1001011001110;
      10'b1100000010:
        _o_sv = 13'b1001011010100;
      10'b1100000011:
        _o_sv = 13'b1001011011010;
      10'b1100000100:
        _o_sv = 13'b1001011100000;
      10'b1100000101:
        _o_sv = 13'b1001011100111;
      10'b1100000110:
        _o_sv = 13'b1001011101101;
      10'b1100000111:
        _o_sv = 13'b1001011110011;
      10'b1100001000:
        _o_sv = 13'b1001011111001;
      10'b1100001001:
        _o_sv = 13'b1001011111111;
      10'b1100001010:
        _o_sv = 13'b1001100000110;
      10'b1100001011:
        _o_sv = 13'b1001100001100;
      10'b1100001100:
        _o_sv = 13'b1001100010010;
      10'b1100001101:
        _o_sv = 13'b1001100011000;
      10'b1100001110:
        _o_sv = 13'b1001100011111;
      10'b1100001111:
        _o_sv = 13'b1001100100101;
      10'b1100010000:
        _o_sv = 13'b1001100101011;
      10'b1100010001:
        _o_sv = 13'b1001100110001;
      10'b1100010010:
        _o_sv = 13'b1001100110111;
      10'b1100010011:
        _o_sv = 13'b1001100111110;
      10'b1100010100:
        _o_sv = 13'b1001101000100;
      10'b1100010101:
        _o_sv = 13'b1001101001010;
      10'b1100010110:
        _o_sv = 13'b1001101010000;
      10'b1100010111:
        _o_sv = 13'b1001101010110;
      10'b1100011000:
        _o_sv = 13'b1001101011101;
      10'b1100011001:
        _o_sv = 13'b1001101100011;
      10'b1100011010:
        _o_sv = 13'b1001101101001;
      10'b1100011011:
        _o_sv = 13'b1001101101111;
      10'b1100011100:
        _o_sv = 13'b1001101110110;
      10'b1100011101:
        _o_sv = 13'b1001101111100;
      10'b1100011110:
        _o_sv = 13'b1001110000010;
      10'b1100011111:
        _o_sv = 13'b1001110001000;
      10'b1100100000:
        _o_sv = 13'b1001110001110;
      10'b1100100001:
        _o_sv = 13'b1001110010101;
      10'b1100100010:
        _o_sv = 13'b1001110011011;
      10'b1100100011:
        _o_sv = 13'b1001110100001;
      10'b1100100100:
        _o_sv = 13'b1001110100111;
      10'b1100100101:
        _o_sv = 13'b1001110101101;
      10'b1100100110:
        _o_sv = 13'b1001110110100;
      10'b1100100111:
        _o_sv = 13'b1001110111010;
      10'b1100101000:
        _o_sv = 13'b1001111000000;
      10'b1100101001:
        _o_sv = 13'b1001111000110;
      10'b1100101010:
        _o_sv = 13'b1001111001100;
      10'b1100101011:
        _o_sv = 13'b1001111010011;
      10'b1100101100:
        _o_sv = 13'b1001111011001;
      10'b1100101101:
        _o_sv = 13'b1001111011111;
      10'b1100101110:
        _o_sv = 13'b1001111100101;
      10'b1100101111:
        _o_sv = 13'b1001111101011;
      10'b1100110000:
        _o_sv = 13'b1001111110010;
      10'b1100110001:
        _o_sv = 13'b1001111111000;
      10'b1100110010:
        _o_sv = 13'b1001111111110;
      10'b1100110011:
        _o_sv = 13'b1010000000100;
      10'b1100110100:
        _o_sv = 13'b1010000001011;
      10'b1100110101:
        _o_sv = 13'b1010000010001;
      10'b1100110110:
        _o_sv = 13'b1010000010111;
      10'b1100110111:
        _o_sv = 13'b1010000011101;
      10'b1100111000:
        _o_sv = 13'b1010000100011;
      10'b1100111001:
        _o_sv = 13'b1010000101010;
      10'b1100111010:
        _o_sv = 13'b1010000110000;
      10'b1100111011:
        _o_sv = 13'b1010000110110;
      10'b1100111100:
        _o_sv = 13'b1010000111100;
      10'b1100111101:
        _o_sv = 13'b1010001000010;
      10'b1100111110:
        _o_sv = 13'b1010001001001;
      10'b1100111111:
        _o_sv = 13'b1010001001111;
      10'b1101000000:
        _o_sv = 13'b1010001010101;
      10'b1101000001:
        _o_sv = 13'b1010001011011;
      10'b1101000010:
        _o_sv = 13'b1010001100001;
      10'b1101000011:
        _o_sv = 13'b1010001101000;
      10'b1101000100:
        _o_sv = 13'b1010001101110;
      10'b1101000101:
        _o_sv = 13'b1010001110100;
      10'b1101000110:
        _o_sv = 13'b1010001111010;
      10'b1101000111:
        _o_sv = 13'b1010010000000;
      10'b1101001000:
        _o_sv = 13'b1010010000111;
      10'b1101001001:
        _o_sv = 13'b1010010001101;
      10'b1101001010:
        _o_sv = 13'b1010010010011;
      10'b1101001011:
        _o_sv = 13'b1010010011001;
      10'b1101001100:
        _o_sv = 13'b1010010011111;
      10'b1101001101:
        _o_sv = 13'b1010010100110;
      10'b1101001110:
        _o_sv = 13'b1010010101100;
      10'b1101001111:
        _o_sv = 13'b1010010110010;
      10'b1101010000:
        _o_sv = 13'b1010010111000;
      10'b1101010001:
        _o_sv = 13'b1010010111110;
      10'b1101010010:
        _o_sv = 13'b1010011000101;
      10'b1101010011:
        _o_sv = 13'b1010011001011;
      10'b1101010100:
        _o_sv = 13'b1010011010001;
      10'b1101010101:
        _o_sv = 13'b1010011010111;
      10'b1101010110:
        _o_sv = 13'b1010011011101;
      10'b1101010111:
        _o_sv = 13'b1010011100100;
      10'b1101011000:
        _o_sv = 13'b1010011101010;
      10'b1101011001:
        _o_sv = 13'b1010011110000;
      10'b1101011010:
        _o_sv = 13'b1010011110110;
      10'b1101011011:
        _o_sv = 13'b1010011111100;
      10'b1101011100:
        _o_sv = 13'b1010100000011;
      10'b1101011101:
        _o_sv = 13'b1010100001001;
      10'b1101011110:
        _o_sv = 13'b1010100001111;
      10'b1101011111:
        _o_sv = 13'b1010100010101;
      10'b1101100000:
        _o_sv = 13'b1010100011011;
      10'b1101100001:
        _o_sv = 13'b1010100100010;
      10'b1101100010:
        _o_sv = 13'b1010100101000;
      10'b1101100011:
        _o_sv = 13'b1010100101110;
      10'b1101100100:
        _o_sv = 13'b1010100110100;
      10'b1101100101:
        _o_sv = 13'b1010100111010;
      10'b1101100110:
        _o_sv = 13'b1010101000001;
      10'b1101100111:
        _o_sv = 13'b1010101000111;
      10'b1101101000:
        _o_sv = 13'b1010101001101;
      10'b1101101001:
        _o_sv = 13'b1010101010011;
      10'b1101101010:
        _o_sv = 13'b1010101011001;
      10'b1101101011:
        _o_sv = 13'b1010101100000;
      10'b1101101100:
        _o_sv = 13'b1010101100110;
      10'b1101101101:
        _o_sv = 13'b1010101101100;
      10'b1101101110:
        _o_sv = 13'b1010101110010;
      10'b1101101111:
        _o_sv = 13'b1010101111000;
      10'b1101110000:
        _o_sv = 13'b1010101111111;
      10'b1101110001:
        _o_sv = 13'b1010110000101;
      10'b1101110010:
        _o_sv = 13'b1010110001011;
      10'b1101110011:
        _o_sv = 13'b1010110010001;
      10'b1101110100:
        _o_sv = 13'b1010110010111;
      10'b1101110101:
        _o_sv = 13'b1010110011101;
      10'b1101110110:
        _o_sv = 13'b1010110100100;
      10'b1101110111:
        _o_sv = 13'b1010110101010;
      10'b1101111000:
        _o_sv = 13'b1010110110000;
      10'b1101111001:
        _o_sv = 13'b1010110110110;
      10'b1101111010:
        _o_sv = 13'b1010110111100;
      10'b1101111011:
        _o_sv = 13'b1010111000011;
      10'b1101111100:
        _o_sv = 13'b1010111001001;
      10'b1101111101:
        _o_sv = 13'b1010111001111;
      10'b1101111110:
        _o_sv = 13'b1010111010101;
      10'b1101111111:
        _o_sv = 13'b1010111011011;
      10'b1110000000:
        _o_sv = 13'b1010111100010;
      10'b1110000001:
        _o_sv = 13'b1010111101000;
      10'b1110000010:
        _o_sv = 13'b1010111101110;
      10'b1110000011:
        _o_sv = 13'b1010111110100;
      10'b1110000100:
        _o_sv = 13'b1010111111010;
      10'b1110000101:
        _o_sv = 13'b1011000000001;
      10'b1110000110:
        _o_sv = 13'b1011000000111;
      10'b1110000111:
        _o_sv = 13'b1011000001101;
      10'b1110001000:
        _o_sv = 13'b1011000010011;
      10'b1110001001:
        _o_sv = 13'b1011000011001;
      10'b1110001010:
        _o_sv = 13'b1011000011111;
      10'b1110001011:
        _o_sv = 13'b1011000100110;
      10'b1110001100:
        _o_sv = 13'b1011000101100;
      10'b1110001101:
        _o_sv = 13'b1011000110010;
      10'b1110001110:
        _o_sv = 13'b1011000111000;
      10'b1110001111:
        _o_sv = 13'b1011000111110;
      10'b1110010000:
        _o_sv = 13'b1011001000101;
      10'b1110010001:
        _o_sv = 13'b1011001001011;
      10'b1110010010:
        _o_sv = 13'b1011001010001;
      10'b1110010011:
        _o_sv = 13'b1011001010111;
      10'b1110010100:
        _o_sv = 13'b1011001011101;
      10'b1110010101:
        _o_sv = 13'b1011001100100;
      10'b1110010110:
        _o_sv = 13'b1011001101010;
      10'b1110010111:
        _o_sv = 13'b1011001110000;
      10'b1110011000:
        _o_sv = 13'b1011001110110;
      10'b1110011001:
        _o_sv = 13'b1011001111100;
      10'b1110011010:
        _o_sv = 13'b1011010000010;
      10'b1110011011:
        _o_sv = 13'b1011010001001;
      10'b1110011100:
        _o_sv = 13'b1011010001111;
      10'b1110011101:
        _o_sv = 13'b1011010010101;
      10'b1110011110:
        _o_sv = 13'b1011010011011;
      10'b1110011111:
        _o_sv = 13'b1011010100001;
      10'b1110100000:
        _o_sv = 13'b1011010101000;
      10'b1110100001:
        _o_sv = 13'b1011010101110;
      10'b1110100010:
        _o_sv = 13'b1011010110100;
      10'b1110100011:
        _o_sv = 13'b1011010111010;
      10'b1110100100:
        _o_sv = 13'b1011011000000;
      10'b1110100101:
        _o_sv = 13'b1011011000110;
      10'b1110100110:
        _o_sv = 13'b1011011001101;
      10'b1110100111:
        _o_sv = 13'b1011011010011;
      10'b1110101000:
        _o_sv = 13'b1011011011001;
      10'b1110101001:
        _o_sv = 13'b1011011011111;
      10'b1110101010:
        _o_sv = 13'b1011011100101;
      10'b1110101011:
        _o_sv = 13'b1011011101100;
      10'b1110101100:
        _o_sv = 13'b1011011110010;
      10'b1110101101:
        _o_sv = 13'b1011011111000;
      10'b1110101110:
        _o_sv = 13'b1011011111110;
      10'b1110101111:
        _o_sv = 13'b1011100000100;
      10'b1110110000:
        _o_sv = 13'b1011100001010;
      10'b1110110001:
        _o_sv = 13'b1011100010001;
      10'b1110110010:
        _o_sv = 13'b1011100010111;
      10'b1110110011:
        _o_sv = 13'b1011100011101;
      10'b1110110100:
        _o_sv = 13'b1011100100011;
      10'b1110110101:
        _o_sv = 13'b1011100101001;
      10'b1110110110:
        _o_sv = 13'b1011100110000;
      10'b1110110111:
        _o_sv = 13'b1011100110110;
      10'b1110111000:
        _o_sv = 13'b1011100111100;
      10'b1110111001:
        _o_sv = 13'b1011101000010;
      10'b1110111010:
        _o_sv = 13'b1011101001000;
      10'b1110111011:
        _o_sv = 13'b1011101001110;
      10'b1110111100:
        _o_sv = 13'b1011101010101;
      10'b1110111101:
        _o_sv = 13'b1011101011011;
      10'b1110111110:
        _o_sv = 13'b1011101100001;
      10'b1110111111:
        _o_sv = 13'b1011101100111;
      10'b1111000000:
        _o_sv = 13'b1011101101101;
      10'b1111000001:
        _o_sv = 13'b1011101110100;
      10'b1111000010:
        _o_sv = 13'b1011101111010;
      10'b1111000011:
        _o_sv = 13'b1011110000000;
      10'b1111000100:
        _o_sv = 13'b1011110000110;
      10'b1111000101:
        _o_sv = 13'b1011110001100;
      10'b1111000110:
        _o_sv = 13'b1011110010010;
      10'b1111000111:
        _o_sv = 13'b1011110011001;
      10'b1111001000:
        _o_sv = 13'b1011110011111;
      10'b1111001001:
        _o_sv = 13'b1011110100101;
      10'b1111001010:
        _o_sv = 13'b1011110101011;
      10'b1111001011:
        _o_sv = 13'b1011110110001;
      10'b1111001100:
        _o_sv = 13'b1011110110111;
      10'b1111001101:
        _o_sv = 13'b1011110111110;
      10'b1111001110:
        _o_sv = 13'b1011111000100;
      10'b1111001111:
        _o_sv = 13'b1011111001010;
      10'b1111010000:
        _o_sv = 13'b1011111010000;
      10'b1111010001:
        _o_sv = 13'b1011111010110;
      10'b1111010010:
        _o_sv = 13'b1011111011101;
      10'b1111010011:
        _o_sv = 13'b1011111100011;
      10'b1111010100:
        _o_sv = 13'b1011111101001;
      10'b1111010101:
        _o_sv = 13'b1011111101111;
      10'b1111010110:
        _o_sv = 13'b1011111110101;
      10'b1111010111:
        _o_sv = 13'b1011111111011;
      10'b1111011000:
        _o_sv = 13'b1100000000010;
      10'b1111011001:
        _o_sv = 13'b1100000001000;
      10'b1111011010:
        _o_sv = 13'b1100000001110;
      10'b1111011011:
        _o_sv = 13'b1100000010100;
      10'b1111011100:
        _o_sv = 13'b1100000011010;
      10'b1111011101:
        _o_sv = 13'b1100000100000;
      10'b1111011110:
        _o_sv = 13'b1100000100111;
      10'b1111011111:
        _o_sv = 13'b1100000101101;
      10'b1111100000:
        _o_sv = 13'b1100000110011;
      10'b1111100001:
        _o_sv = 13'b1100000111001;
      10'b1111100010:
        _o_sv = 13'b1100000111111;
      10'b1111100011:
        _o_sv = 13'b1100001000101;
      10'b1111100100:
        _o_sv = 13'b1100001001100;
      10'b1111100101:
        _o_sv = 13'b1100001010010;
      10'b1111100110:
        _o_sv = 13'b1100001011000;
      10'b1111100111:
        _o_sv = 13'b1100001011110;
      10'b1111101000:
        _o_sv = 13'b1100001100100;
      10'b1111101001:
        _o_sv = 13'b1100001101010;
      10'b1111101010:
        _o_sv = 13'b1100001110001;
      10'b1111101011:
        _o_sv = 13'b1100001110111;
      10'b1111101100:
        _o_sv = 13'b1100001111101;
      10'b1111101101:
        _o_sv = 13'b1100010000011;
      10'b1111101110:
        _o_sv = 13'b1100010001001;
      10'b1111101111:
        _o_sv = 13'b1100010001111;
      10'b1111110000:
        _o_sv = 13'b1100010010110;
      10'b1111110001:
        _o_sv = 13'b1100010011100;
      10'b1111110010:
        _o_sv = 13'b1100010100010;
      10'b1111110011:
        _o_sv = 13'b1100010101000;
      10'b1111110100:
        _o_sv = 13'b1100010101110;
      10'b1111110101:
        _o_sv = 13'b1100010110100;
      10'b1111110110:
        _o_sv = 13'b1100010111011;
      10'b1111110111:
        _o_sv = 13'b1100011000001;
      10'b1111111000:
        _o_sv = 13'b1100011000111;
      10'b1111111001:
        _o_sv = 13'b1100011001101;
      10'b1111111010:
        _o_sv = 13'b1100011010011;
      10'b1111111011:
        _o_sv = 13'b1100011011001;
      10'b1111111100:
        _o_sv = 13'b1100011100000;
      10'b1111111101:
        _o_sv = 13'b1100011100110;
      10'b1111111110:
        _o_sv = 13'b1100011101100;
      10'b1111111111:
        _o_sv = 13'b1100011110010;
      11'b10000000000:
        _o_sv = 13'b1100011111000;
      11'b10000000001:
        _o_sv = 13'b1100011111110;
      11'b10000000010:
        _o_sv = 13'b1100100000101;
      11'b10000000011:
        _o_sv = 13'b1100100001011;
      11'b10000000100:
        _o_sv = 13'b1100100010001;
      11'b10000000101:
        _o_sv = 13'b1100100010111;
      11'b10000000110:
        _o_sv = 13'b1100100011101;
      11'b10000000111:
        _o_sv = 13'b1100100100011;
      11'b10000001000:
        _o_sv = 13'b1100100101010;
      11'b10000001001:
        _o_sv = 13'b1100100110000;
      11'b10000001010:
        _o_sv = 13'b1100100110110;
      11'b10000001011:
        _o_sv = 13'b1100100111100;
      11'b10000001100:
        _o_sv = 13'b1100101000010;
      11'b10000001101:
        _o_sv = 13'b1100101001000;
      11'b10000001110:
        _o_sv = 13'b1100101001110;
      11'b10000001111:
        _o_sv = 13'b1100101010101;
      11'b10000010000:
        _o_sv = 13'b1100101011011;
      11'b10000010001:
        _o_sv = 13'b1100101100001;
      11'b10000010010:
        _o_sv = 13'b1100101100111;
      11'b10000010011:
        _o_sv = 13'b1100101101101;
      11'b10000010100:
        _o_sv = 13'b1100101110011;
      11'b10000010101:
        _o_sv = 13'b1100101111010;
      11'b10000010110:
        _o_sv = 13'b1100110000000;
      11'b10000010111:
        _o_sv = 13'b1100110000110;
      11'b10000011000:
        _o_sv = 13'b1100110001100;
      11'b10000011001:
        _o_sv = 13'b1100110010010;
      11'b10000011010:
        _o_sv = 13'b1100110011000;
      11'b10000011011:
        _o_sv = 13'b1100110011111;
      11'b10000011100:
        _o_sv = 13'b1100110100101;
      11'b10000011101:
        _o_sv = 13'b1100110101011;
      11'b10000011110:
        _o_sv = 13'b1100110110001;
      11'b10000011111:
        _o_sv = 13'b1100110110111;
      11'b10000100000:
        _o_sv = 13'b1100110111101;
      11'b10000100001:
        _o_sv = 13'b1100111000011;
      11'b10000100010:
        _o_sv = 13'b1100111001010;
      11'b10000100011:
        _o_sv = 13'b1100111010000;
      11'b10000100100:
        _o_sv = 13'b1100111010110;
      11'b10000100101:
        _o_sv = 13'b1100111011100;
      11'b10000100110:
        _o_sv = 13'b1100111100010;
      11'b10000100111:
        _o_sv = 13'b1100111101000;
      11'b10000101000:
        _o_sv = 13'b1100111101111;
      11'b10000101001:
        _o_sv = 13'b1100111110101;
      11'b10000101010:
        _o_sv = 13'b1100111111011;
      11'b10000101011:
        _o_sv = 13'b1101000000001;
      11'b10000101100:
        _o_sv = 13'b1101000000111;
      11'b10000101101:
        _o_sv = 13'b1101000001101;
      11'b10000101110:
        _o_sv = 13'b1101000010011;
      11'b10000101111:
        _o_sv = 13'b1101000011010;
      11'b10000110000:
        _o_sv = 13'b1101000100000;
      11'b10000110001:
        _o_sv = 13'b1101000100110;
      11'b10000110010:
        _o_sv = 13'b1101000101100;
      11'b10000110011:
        _o_sv = 13'b1101000110010;
      11'b10000110100:
        _o_sv = 13'b1101000111000;
      11'b10000110101:
        _o_sv = 13'b1101000111110;
      11'b10000110110:
        _o_sv = 13'b1101001000101;
      11'b10000110111:
        _o_sv = 13'b1101001001011;
      11'b10000111000:
        _o_sv = 13'b1101001010001;
      11'b10000111001:
        _o_sv = 13'b1101001010111;
      11'b10000111010:
        _o_sv = 13'b1101001011101;
      11'b10000111011:
        _o_sv = 13'b1101001100011;
      11'b10000111100:
        _o_sv = 13'b1101001101010;
      11'b10000111101:
        _o_sv = 13'b1101001110000;
      11'b10000111110:
        _o_sv = 13'b1101001110110;
      11'b10000111111:
        _o_sv = 13'b1101001111100;
      11'b10001000000:
        _o_sv = 13'b1101010000010;
      11'b10001000001:
        _o_sv = 13'b1101010001000;
      11'b10001000010:
        _o_sv = 13'b1101010001110;
      11'b10001000011:
        _o_sv = 13'b1101010010101;
      11'b10001000100:
        _o_sv = 13'b1101010011011;
      11'b10001000101:
        _o_sv = 13'b1101010100001;
      11'b10001000110:
        _o_sv = 13'b1101010100111;
      11'b10001000111:
        _o_sv = 13'b1101010101101;
      11'b10001001000:
        _o_sv = 13'b1101010110011;
      11'b10001001001:
        _o_sv = 13'b1101010111001;
      11'b10001001010:
        _o_sv = 13'b1101011000000;
      11'b10001001011:
        _o_sv = 13'b1101011000110;
      11'b10001001100:
        _o_sv = 13'b1101011001100;
      11'b10001001101:
        _o_sv = 13'b1101011010010;
      11'b10001001110:
        _o_sv = 13'b1101011011000;
      11'b10001001111:
        _o_sv = 13'b1101011011110;
      11'b10001010000:
        _o_sv = 13'b1101011100100;
      11'b10001010001:
        _o_sv = 13'b1101011101011;
      11'b10001010010:
        _o_sv = 13'b1101011110001;
      11'b10001010011:
        _o_sv = 13'b1101011110111;
      11'b10001010100:
        _o_sv = 13'b1101011111101;
      11'b10001010101:
        _o_sv = 13'b1101100000011;
      11'b10001010110:
        _o_sv = 13'b1101100001001;
      11'b10001010111:
        _o_sv = 13'b1101100001111;
      11'b10001011000:
        _o_sv = 13'b1101100010110;
      11'b10001011001:
        _o_sv = 13'b1101100011100;
      11'b10001011010:
        _o_sv = 13'b1101100100010;
      11'b10001011011:
        _o_sv = 13'b1101100101000;
      11'b10001011100:
        _o_sv = 13'b1101100101110;
      11'b10001011101:
        _o_sv = 13'b1101100110100;
      11'b10001011110:
        _o_sv = 13'b1101100111010;
      11'b10001011111:
        _o_sv = 13'b1101101000001;
      11'b10001100000:
        _o_sv = 13'b1101101000111;
      11'b10001100001:
        _o_sv = 13'b1101101001101;
      11'b10001100010:
        _o_sv = 13'b1101101010011;
      11'b10001100011:
        _o_sv = 13'b1101101011001;
      11'b10001100100:
        _o_sv = 13'b1101101011111;
      11'b10001100101:
        _o_sv = 13'b1101101100101;
      11'b10001100110:
        _o_sv = 13'b1101101101100;
      11'b10001100111:
        _o_sv = 13'b1101101110010;
      11'b10001101000:
        _o_sv = 13'b1101101111000;
      11'b10001101001:
        _o_sv = 13'b1101101111110;
      11'b10001101010:
        _o_sv = 13'b1101110000100;
      11'b10001101011:
        _o_sv = 13'b1101110001010;
      11'b10001101100:
        _o_sv = 13'b1101110010000;
      11'b10001101101:
        _o_sv = 13'b1101110010110;
      11'b10001101110:
        _o_sv = 13'b1101110011101;
      11'b10001101111:
        _o_sv = 13'b1101110100011;
      11'b10001110000:
        _o_sv = 13'b1101110101001;
      11'b10001110001:
        _o_sv = 13'b1101110101111;
      11'b10001110010:
        _o_sv = 13'b1101110110101;
      11'b10001110011:
        _o_sv = 13'b1101110111011;
      11'b10001110100:
        _o_sv = 13'b1101111000001;
      11'b10001110101:
        _o_sv = 13'b1101111001000;
      11'b10001110110:
        _o_sv = 13'b1101111001110;
      11'b10001110111:
        _o_sv = 13'b1101111010100;
      11'b10001111000:
        _o_sv = 13'b1101111011010;
      11'b10001111001:
        _o_sv = 13'b1101111100000;
      11'b10001111010:
        _o_sv = 13'b1101111100110;
      11'b10001111011:
        _o_sv = 13'b1101111101100;
      11'b10001111100:
        _o_sv = 13'b1101111110010;
      11'b10001111101:
        _o_sv = 13'b1101111111001;
      11'b10001111110:
        _o_sv = 13'b1101111111111;
      11'b10001111111:
        _o_sv = 13'b1110000000101;
      11'b10010000000:
        _o_sv = 13'b1110000001011;
      11'b10010000001:
        _o_sv = 13'b1110000010001;
      11'b10010000010:
        _o_sv = 13'b1110000010111;
      11'b10010000011:
        _o_sv = 13'b1110000011101;
      11'b10010000100:
        _o_sv = 13'b1110000100100;
      11'b10010000101:
        _o_sv = 13'b1110000101010;
      11'b10010000110:
        _o_sv = 13'b1110000110000;
      11'b10010000111:
        _o_sv = 13'b1110000110110;
      11'b10010001000:
        _o_sv = 13'b1110000111100;
      11'b10010001001:
        _o_sv = 13'b1110001000010;
      11'b10010001010:
        _o_sv = 13'b1110001001000;
      11'b10010001011:
        _o_sv = 13'b1110001001110;
      11'b10010001100:
        _o_sv = 13'b1110001010101;
      11'b10010001101:
        _o_sv = 13'b1110001011011;
      11'b10010001110:
        _o_sv = 13'b1110001100001;
      11'b10010001111:
        _o_sv = 13'b1110001100111;
      11'b10010010000:
        _o_sv = 13'b1110001101101;
      11'b10010010001:
        _o_sv = 13'b1110001110011;
      11'b10010010010:
        _o_sv = 13'b1110001111001;
      11'b10010010011:
        _o_sv = 13'b1110001111111;
      11'b10010010100:
        _o_sv = 13'b1110010000110;
      11'b10010010101:
        _o_sv = 13'b1110010001100;
      11'b10010010110:
        _o_sv = 13'b1110010010010;
      11'b10010010111:
        _o_sv = 13'b1110010011000;
      11'b10010011000:
        _o_sv = 13'b1110010011110;
      11'b10010011001:
        _o_sv = 13'b1110010100100;
      11'b10010011010:
        _o_sv = 13'b1110010101010;
      11'b10010011011:
        _o_sv = 13'b1110010110000;
      11'b10010011100:
        _o_sv = 13'b1110010110111;
      11'b10010011101:
        _o_sv = 13'b1110010111101;
      11'b10010011110:
        _o_sv = 13'b1110011000011;
      11'b10010011111:
        _o_sv = 13'b1110011001001;
      11'b10010100000:
        _o_sv = 13'b1110011001111;
      11'b10010100001:
        _o_sv = 13'b1110011010101;
      11'b10010100010:
        _o_sv = 13'b1110011011011;
      11'b10010100011:
        _o_sv = 13'b1110011100001;
      11'b10010100100:
        _o_sv = 13'b1110011101000;
      11'b10010100101:
        _o_sv = 13'b1110011101110;
      11'b10010100110:
        _o_sv = 13'b1110011110100;
      11'b10010100111:
        _o_sv = 13'b1110011111010;
      11'b10010101000:
        _o_sv = 13'b1110100000000;
      11'b10010101001:
        _o_sv = 13'b1110100000110;
      11'b10010101010:
        _o_sv = 13'b1110100001100;
      11'b10010101011:
        _o_sv = 13'b1110100010010;
      11'b10010101100:
        _o_sv = 13'b1110100011000;
      11'b10010101101:
        _o_sv = 13'b1110100011111;
      11'b10010101110:
        _o_sv = 13'b1110100100101;
      11'b10010101111:
        _o_sv = 13'b1110100101011;
      11'b10010110000:
        _o_sv = 13'b1110100110001;
      11'b10010110001:
        _o_sv = 13'b1110100110111;
      11'b10010110010:
        _o_sv = 13'b1110100111101;
      11'b10010110011:
        _o_sv = 13'b1110101000011;
      11'b10010110100:
        _o_sv = 13'b1110101001001;
      11'b10010110101:
        _o_sv = 13'b1110101010000;
      11'b10010110110:
        _o_sv = 13'b1110101010110;
      11'b10010110111:
        _o_sv = 13'b1110101011100;
      11'b10010111000:
        _o_sv = 13'b1110101100010;
      11'b10010111001:
        _o_sv = 13'b1110101101000;
      11'b10010111010:
        _o_sv = 13'b1110101101110;
      11'b10010111011:
        _o_sv = 13'b1110101110100;
      11'b10010111100:
        _o_sv = 13'b1110101111010;
      11'b10010111101:
        _o_sv = 13'b1110110000000;
      11'b10010111110:
        _o_sv = 13'b1110110000111;
      11'b10010111111:
        _o_sv = 13'b1110110001101;
      11'b10011000000:
        _o_sv = 13'b1110110010011;
      11'b10011000001:
        _o_sv = 13'b1110110011001;
      11'b10011000010:
        _o_sv = 13'b1110110011111;
      11'b10011000011:
        _o_sv = 13'b1110110100101;
      11'b10011000100:
        _o_sv = 13'b1110110101011;
      11'b10011000101:
        _o_sv = 13'b1110110110001;
      11'b10011000110:
        _o_sv = 13'b1110110110111;
      11'b10011000111:
        _o_sv = 13'b1110110111110;
      11'b10011001000:
        _o_sv = 13'b1110111000100;
      11'b10011001001:
        _o_sv = 13'b1110111001010;
      11'b10011001010:
        _o_sv = 13'b1110111010000;
      11'b10011001011:
        _o_sv = 13'b1110111010110;
      11'b10011001100:
        _o_sv = 13'b1110111011100;
      11'b10011001101:
        _o_sv = 13'b1110111100010;
      11'b10011001110:
        _o_sv = 13'b1110111101000;
      11'b10011001111:
        _o_sv = 13'b1110111101110;
      11'b10011010000:
        _o_sv = 13'b1110111110101;
      11'b10011010001:
        _o_sv = 13'b1110111111011;
      11'b10011010010:
        _o_sv = 13'b1111000000001;
      11'b10011010011:
        _o_sv = 13'b1111000000111;
      11'b10011010100:
        _o_sv = 13'b1111000001101;
      11'b10011010101:
        _o_sv = 13'b1111000010011;
      11'b10011010110:
        _o_sv = 13'b1111000011001;
      11'b10011010111:
        _o_sv = 13'b1111000011111;
      11'b10011011000:
        _o_sv = 13'b1111000100101;
      11'b10011011001:
        _o_sv = 13'b1111000101100;
      11'b10011011010:
        _o_sv = 13'b1111000110010;
      11'b10011011011:
        _o_sv = 13'b1111000111000;
      11'b10011011100:
        _o_sv = 13'b1111000111110;
      11'b10011011101:
        _o_sv = 13'b1111001000100;
      11'b10011011110:
        _o_sv = 13'b1111001001010;
      11'b10011011111:
        _o_sv = 13'b1111001010000;
      11'b10011100000:
        _o_sv = 13'b1111001010110;
      11'b10011100001:
        _o_sv = 13'b1111001011100;
      11'b10011100010:
        _o_sv = 13'b1111001100010;
      11'b10011100011:
        _o_sv = 13'b1111001101001;
      11'b10011100100:
        _o_sv = 13'b1111001101111;
      11'b10011100101:
        _o_sv = 13'b1111001110101;
      11'b10011100110:
        _o_sv = 13'b1111001111011;
      11'b10011100111:
        _o_sv = 13'b1111010000001;
      11'b10011101000:
        _o_sv = 13'b1111010000111;
      11'b10011101001:
        _o_sv = 13'b1111010001101;
      11'b10011101010:
        _o_sv = 13'b1111010010011;
      11'b10011101011:
        _o_sv = 13'b1111010011001;
      11'b10011101100:
        _o_sv = 13'b1111010100000;
      11'b10011101101:
        _o_sv = 13'b1111010100110;
      11'b10011101110:
        _o_sv = 13'b1111010101100;
      11'b10011101111:
        _o_sv = 13'b1111010110010;
      11'b10011110000:
        _o_sv = 13'b1111010111000;
      11'b10011110001:
        _o_sv = 13'b1111010111110;
      11'b10011110010:
        _o_sv = 13'b1111011000100;
      11'b10011110011:
        _o_sv = 13'b1111011001010;
      11'b10011110100:
        _o_sv = 13'b1111011010000;
      11'b10011110101:
        _o_sv = 13'b1111011010110;
      11'b10011110110:
        _o_sv = 13'b1111011011101;
      11'b10011110111:
        _o_sv = 13'b1111011100011;
      11'b10011111000:
        _o_sv = 13'b1111011101001;
      11'b10011111001:
        _o_sv = 13'b1111011101111;
      11'b10011111010:
        _o_sv = 13'b1111011110101;
      11'b10011111011:
        _o_sv = 13'b1111011111011;
      11'b10011111100:
        _o_sv = 13'b1111100000001;
      11'b10011111101:
        _o_sv = 13'b1111100000111;
      11'b10011111110:
        _o_sv = 13'b1111100001101;
      11'b10011111111:
        _o_sv = 13'b1111100010011;
      11'b10100000000:
        _o_sv = 13'b1111100011001;
      11'b10100000001:
        _o_sv = 13'b1111100100000;
      11'b10100000010:
        _o_sv = 13'b1111100100110;
      11'b10100000011:
        _o_sv = 13'b1111100101100;
      11'b10100000100:
        _o_sv = 13'b1111100110010;
      11'b10100000101:
        _o_sv = 13'b1111100111000;
      11'b10100000110:
        _o_sv = 13'b1111100111110;
      11'b10100000111:
        _o_sv = 13'b1111101000100;
      11'b10100001000:
        _o_sv = 13'b1111101001010;
      11'b10100001001:
        _o_sv = 13'b1111101010000;
      11'b10100001010:
        _o_sv = 13'b1111101010110;
      11'b10100001011:
        _o_sv = 13'b1111101011101;
      11'b10100001100:
        _o_sv = 13'b1111101100011;
      11'b10100001101:
        _o_sv = 13'b1111101101001;
      11'b10100001110:
        _o_sv = 13'b1111101101111;
      11'b10100001111:
        _o_sv = 13'b1111101110101;
      11'b10100010000:
        _o_sv = 13'b1111101111011;
      11'b10100010001:
        _o_sv = 13'b1111110000001;
      11'b10100010010:
        _o_sv = 13'b1111110000111;
      11'b10100010011:
        _o_sv = 13'b1111110001101;
      11'b10100010100:
        _o_sv = 13'b1111110010011;
      11'b10100010101:
        _o_sv = 13'b1111110011001;
      11'b10100010110:
        _o_sv = 13'b1111110011111;
      11'b10100010111:
        _o_sv = 13'b1111110100110;
      11'b10100011000:
        _o_sv = 13'b1111110101100;
      11'b10100011001:
        _o_sv = 13'b1111110110010;
      11'b10100011010:
        _o_sv = 13'b1111110111000;
      11'b10100011011:
        _o_sv = 13'b1111110111110;
      11'b10100011100:
        _o_sv = 13'b1111111000100;
      11'b10100011101:
        _o_sv = 13'b1111111001010;
      11'b10100011110:
        _o_sv = 13'b1111111010000;
      11'b10100011111:
        _o_sv = 13'b1111111010110;
      11'b10100100000:
        _o_sv = 13'b1111111011100;
      11'b10100100001:
        _o_sv = 13'b1111111100010;
      11'b10100100010:
        _o_sv = 13'b1111111101001;
      11'b10100100011:
        _o_sv = 13'b1111111101111;
      11'b10100100100:
        _o_sv = 13'b1111111110101;
      11'b10100100101:
        _o_sv = 13'b1111111111011;
      11'b10100100110:
        _o_sv = 14'b10000000000001;
      11'b10100100111:
        _o_sv = 14'b10000000000111;
      11'b10100101000:
        _o_sv = 14'b10000000001101;
      11'b10100101001:
        _o_sv = 14'b10000000010011;
      11'b10100101010:
        _o_sv = 14'b10000000011001;
      11'b10100101011:
        _o_sv = 14'b10000000011111;
      11'b10100101100:
        _o_sv = 14'b10000000100101;
      11'b10100101101:
        _o_sv = 14'b10000000101011;
      11'b10100101110:
        _o_sv = 14'b10000000110010;
      11'b10100101111:
        _o_sv = 14'b10000000111000;
      11'b10100110000:
        _o_sv = 14'b10000000111110;
      11'b10100110001:
        _o_sv = 14'b10000001000100;
      11'b10100110010:
        _o_sv = 14'b10000001001010;
      11'b10100110011:
        _o_sv = 14'b10000001010000;
      11'b10100110100:
        _o_sv = 14'b10000001010110;
      11'b10100110101:
        _o_sv = 14'b10000001011100;
      11'b10100110110:
        _o_sv = 14'b10000001100010;
      11'b10100110111:
        _o_sv = 14'b10000001101000;
      11'b10100111000:
        _o_sv = 14'b10000001101110;
      11'b10100111001:
        _o_sv = 14'b10000001110100;
      11'b10100111010:
        _o_sv = 14'b10000001111010;
      11'b10100111011:
        _o_sv = 14'b10000010000001;
      11'b10100111100:
        _o_sv = 14'b10000010000111;
      11'b10100111101:
        _o_sv = 14'b10000010001101;
      11'b10100111110:
        _o_sv = 14'b10000010010011;
      11'b10100111111:
        _o_sv = 14'b10000010011001;
      11'b10101000000:
        _o_sv = 14'b10000010011111;
      11'b10101000001:
        _o_sv = 14'b10000010100101;
      11'b10101000010:
        _o_sv = 14'b10000010101011;
      11'b10101000011:
        _o_sv = 14'b10000010110001;
      11'b10101000100:
        _o_sv = 14'b10000010110111;
      11'b10101000101:
        _o_sv = 14'b10000010111101;
      11'b10101000110:
        _o_sv = 14'b10000011000011;
      11'b10101000111:
        _o_sv = 14'b10000011001001;
      11'b10101001000:
        _o_sv = 14'b10000011010000;
      11'b10101001001:
        _o_sv = 14'b10000011010110;
      11'b10101001010:
        _o_sv = 14'b10000011011100;
      11'b10101001011:
        _o_sv = 14'b10000011100010;
      11'b10101001100:
        _o_sv = 14'b10000011101000;
      11'b10101001101:
        _o_sv = 14'b10000011101110;
      11'b10101001110:
        _o_sv = 14'b10000011110100;
      11'b10101001111:
        _o_sv = 14'b10000011111010;
      11'b10101010000:
        _o_sv = 14'b10000100000000;
      11'b10101010001:
        _o_sv = 14'b10000100000110;
      11'b10101010010:
        _o_sv = 14'b10000100001100;
      11'b10101010011:
        _o_sv = 14'b10000100010010;
      11'b10101010100:
        _o_sv = 14'b10000100011000;
      11'b10101010101:
        _o_sv = 14'b10000100011110;
      11'b10101010110:
        _o_sv = 14'b10000100100101;
      11'b10101010111:
        _o_sv = 14'b10000100101011;
      11'b10101011000:
        _o_sv = 14'b10000100110001;
      11'b10101011001:
        _o_sv = 14'b10000100110111;
      11'b10101011010:
        _o_sv = 14'b10000100111101;
      11'b10101011011:
        _o_sv = 14'b10000101000011;
      11'b10101011100:
        _o_sv = 14'b10000101001001;
      11'b10101011101:
        _o_sv = 14'b10000101001111;
      11'b10101011110:
        _o_sv = 14'b10000101010101;
      11'b10101011111:
        _o_sv = 14'b10000101011011;
      11'b10101100000:
        _o_sv = 14'b10000101100001;
      11'b10101100001:
        _o_sv = 14'b10000101100111;
      11'b10101100010:
        _o_sv = 14'b10000101101101;
      11'b10101100011:
        _o_sv = 14'b10000101110011;
      11'b10101100100:
        _o_sv = 14'b10000101111001;
      11'b10101100101:
        _o_sv = 14'b10000110000000;
      11'b10101100110:
        _o_sv = 14'b10000110000110;
      11'b10101100111:
        _o_sv = 14'b10000110001100;
      11'b10101101000:
        _o_sv = 14'b10000110010010;
      11'b10101101001:
        _o_sv = 14'b10000110011000;
      11'b10101101010:
        _o_sv = 14'b10000110011110;
      11'b10101101011:
        _o_sv = 14'b10000110100100;
      11'b10101101100:
        _o_sv = 14'b10000110101010;
      11'b10101101101:
        _o_sv = 14'b10000110110000;
      11'b10101101110:
        _o_sv = 14'b10000110110110;
      11'b10101101111:
        _o_sv = 14'b10000110111100;
      11'b10101110000:
        _o_sv = 14'b10000111000010;
      11'b10101110001:
        _o_sv = 14'b10000111001000;
      11'b10101110010:
        _o_sv = 14'b10000111001110;
      11'b10101110011:
        _o_sv = 14'b10000111010100;
      11'b10101110100:
        _o_sv = 14'b10000111011010;
      11'b10101110101:
        _o_sv = 14'b10000111100001;
      11'b10101110110:
        _o_sv = 14'b10000111100111;
      11'b10101110111:
        _o_sv = 14'b10000111101101;
      11'b10101111000:
        _o_sv = 14'b10000111110011;
      11'b10101111001:
        _o_sv = 14'b10000111111001;
      11'b10101111010:
        _o_sv = 14'b10000111111111;
      11'b10101111011:
        _o_sv = 14'b10001000000101;
      11'b10101111100:
        _o_sv = 14'b10001000001011;
      11'b10101111101:
        _o_sv = 14'b10001000010001;
      11'b10101111110:
        _o_sv = 14'b10001000010111;
      11'b10101111111:
        _o_sv = 14'b10001000011101;
      11'b10110000000:
        _o_sv = 14'b10001000100011;
      11'b10110000001:
        _o_sv = 14'b10001000101001;
      11'b10110000010:
        _o_sv = 14'b10001000101111;
      11'b10110000011:
        _o_sv = 14'b10001000110101;
      11'b10110000100:
        _o_sv = 14'b10001000111011;
      11'b10110000101:
        _o_sv = 14'b10001001000001;
      11'b10110000110:
        _o_sv = 14'b10001001000111;
      11'b10110000111:
        _o_sv = 14'b10001001001110;
      11'b10110001000:
        _o_sv = 14'b10001001010100;
      11'b10110001001:
        _o_sv = 14'b10001001011010;
      11'b10110001010:
        _o_sv = 14'b10001001100000;
      11'b10110001011:
        _o_sv = 14'b10001001100110;
      11'b10110001100:
        _o_sv = 14'b10001001101100;
      11'b10110001101:
        _o_sv = 14'b10001001110010;
      11'b10110001110:
        _o_sv = 14'b10001001111000;
      11'b10110001111:
        _o_sv = 14'b10001001111110;
      11'b10110010000:
        _o_sv = 14'b10001010000100;
      11'b10110010001:
        _o_sv = 14'b10001010001010;
      11'b10110010010:
        _o_sv = 14'b10001010010000;
      11'b10110010011:
        _o_sv = 14'b10001010010110;
      11'b10110010100:
        _o_sv = 14'b10001010011100;
      11'b10110010101:
        _o_sv = 14'b10001010100010;
      11'b10110010110:
        _o_sv = 14'b10001010101000;
      11'b10110010111:
        _o_sv = 14'b10001010101110;
      11'b10110011000:
        _o_sv = 14'b10001010110100;
      11'b10110011001:
        _o_sv = 14'b10001010111010;
      11'b10110011010:
        _o_sv = 14'b10001011000000;
      11'b10110011011:
        _o_sv = 14'b10001011000111;
      11'b10110011100:
        _o_sv = 14'b10001011001101;
      11'b10110011101:
        _o_sv = 14'b10001011010011;
      11'b10110011110:
        _o_sv = 14'b10001011011001;
      11'b10110011111:
        _o_sv = 14'b10001011011111;
      11'b10110100000:
        _o_sv = 14'b10001011100101;
      11'b10110100001:
        _o_sv = 14'b10001011101011;
      11'b10110100010:
        _o_sv = 14'b10001011110001;
      11'b10110100011:
        _o_sv = 14'b10001011110111;
      11'b10110100100:
        _o_sv = 14'b10001011111101;
      11'b10110100101:
        _o_sv = 14'b10001100000011;
      11'b10110100110:
        _o_sv = 14'b10001100001001;
      11'b10110100111:
        _o_sv = 14'b10001100001111;
      11'b10110101000:
        _o_sv = 14'b10001100010101;
      11'b10110101001:
        _o_sv = 14'b10001100011011;
      11'b10110101010:
        _o_sv = 14'b10001100100001;
      11'b10110101011:
        _o_sv = 14'b10001100100111;
      11'b10110101100:
        _o_sv = 14'b10001100101101;
      11'b10110101101:
        _o_sv = 14'b10001100110011;
      11'b10110101110:
        _o_sv = 14'b10001100111001;
      11'b10110101111:
        _o_sv = 14'b10001100111111;
      11'b10110110000:
        _o_sv = 14'b10001101000101;
      11'b10110110001:
        _o_sv = 14'b10001101001011;
      11'b10110110010:
        _o_sv = 14'b10001101010010;
      11'b10110110011:
        _o_sv = 14'b10001101011000;
      11'b10110110100:
        _o_sv = 14'b10001101011110;
      11'b10110110101:
        _o_sv = 14'b10001101100100;
      11'b10110110110:
        _o_sv = 14'b10001101101010;
      11'b10110110111:
        _o_sv = 14'b10001101110000;
      11'b10110111000:
        _o_sv = 14'b10001101110110;
      11'b10110111001:
        _o_sv = 14'b10001101111100;
      11'b10110111010:
        _o_sv = 14'b10001110000010;
      11'b10110111011:
        _o_sv = 14'b10001110001000;
      11'b10110111100:
        _o_sv = 14'b10001110001110;
      11'b10110111101:
        _o_sv = 14'b10001110010100;
      11'b10110111110:
        _o_sv = 14'b10001110011010;
      11'b10110111111:
        _o_sv = 14'b10001110100000;
      11'b10111000000:
        _o_sv = 14'b10001110100110;
      11'b10111000001:
        _o_sv = 14'b10001110101100;
      11'b10111000010:
        _o_sv = 14'b10001110110010;
      11'b10111000011:
        _o_sv = 14'b10001110111000;
      11'b10111000100:
        _o_sv = 14'b10001110111110;
      11'b10111000101:
        _o_sv = 14'b10001111000100;
      11'b10111000110:
        _o_sv = 14'b10001111001010;
      11'b10111000111:
        _o_sv = 14'b10001111010000;
      11'b10111001000:
        _o_sv = 14'b10001111010110;
      11'b10111001001:
        _o_sv = 14'b10001111011100;
      11'b10111001010:
        _o_sv = 14'b10001111100010;
      11'b10111001011:
        _o_sv = 14'b10001111101000;
      11'b10111001100:
        _o_sv = 14'b10001111101110;
      11'b10111001101:
        _o_sv = 14'b10001111110100;
      11'b10111001110:
        _o_sv = 14'b10001111111010;
      11'b10111001111:
        _o_sv = 14'b10010000000001;
      11'b10111010000:
        _o_sv = 14'b10010000000111;
      11'b10111010001:
        _o_sv = 14'b10010000001101;
      11'b10111010010:
        _o_sv = 14'b10010000010011;
      11'b10111010011:
        _o_sv = 14'b10010000011001;
      11'b10111010100:
        _o_sv = 14'b10010000011111;
      11'b10111010101:
        _o_sv = 14'b10010000100101;
      11'b10111010110:
        _o_sv = 14'b10010000101011;
      11'b10111010111:
        _o_sv = 14'b10010000110001;
      11'b10111011000:
        _o_sv = 14'b10010000110111;
      11'b10111011001:
        _o_sv = 14'b10010000111101;
      11'b10111011010:
        _o_sv = 14'b10010001000011;
      11'b10111011011:
        _o_sv = 14'b10010001001001;
      11'b10111011100:
        _o_sv = 14'b10010001001111;
      11'b10111011101:
        _o_sv = 14'b10010001010101;
      11'b10111011110:
        _o_sv = 14'b10010001011011;
      11'b10111011111:
        _o_sv = 14'b10010001100001;
      11'b10111100000:
        _o_sv = 14'b10010001100111;
      11'b10111100001:
        _o_sv = 14'b10010001101101;
      11'b10111100010:
        _o_sv = 14'b10010001110011;
      11'b10111100011:
        _o_sv = 14'b10010001111001;
      11'b10111100100:
        _o_sv = 14'b10010001111111;
      11'b10111100101:
        _o_sv = 14'b10010010000101;
      11'b10111100110:
        _o_sv = 14'b10010010001011;
      11'b10111100111:
        _o_sv = 14'b10010010010001;
      11'b10111101000:
        _o_sv = 14'b10010010010111;
      11'b10111101001:
        _o_sv = 14'b10010010011101;
      11'b10111101010:
        _o_sv = 14'b10010010100011;
      11'b10111101011:
        _o_sv = 14'b10010010101001;
      11'b10111101100:
        _o_sv = 14'b10010010101111;
      11'b10111101101:
        _o_sv = 14'b10010010110101;
      11'b10111101110:
        _o_sv = 14'b10010010111011;
      11'b10111101111:
        _o_sv = 14'b10010011000001;
      11'b10111110000:
        _o_sv = 14'b10010011000111;
      11'b10111110001:
        _o_sv = 14'b10010011001101;
      11'b10111110010:
        _o_sv = 14'b10010011010011;
      11'b10111110011:
        _o_sv = 14'b10010011011001;
      11'b10111110100:
        _o_sv = 14'b10010011011111;
      11'b10111110101:
        _o_sv = 14'b10010011100101;
      11'b10111110110:
        _o_sv = 14'b10010011101011;
      11'b10111110111:
        _o_sv = 14'b10010011110001;
      11'b10111111000:
        _o_sv = 14'b10010011110111;
      11'b10111111001:
        _o_sv = 14'b10010011111101;
      11'b10111111010:
        _o_sv = 14'b10010100000011;
      11'b10111111011:
        _o_sv = 14'b10010100001001;
      11'b10111111100:
        _o_sv = 14'b10010100001111;
      11'b10111111101:
        _o_sv = 14'b10010100010110;
      11'b10111111110:
        _o_sv = 14'b10010100011100;
      11'b10111111111:
        _o_sv = 14'b10010100100010;
      11'b11000000000:
        _o_sv = 14'b10010100101000;
      11'b11000000001:
        _o_sv = 14'b10010100101110;
      11'b11000000010:
        _o_sv = 14'b10010100110100;
      11'b11000000011:
        _o_sv = 14'b10010100111010;
      11'b11000000100:
        _o_sv = 14'b10010101000000;
      11'b11000000101:
        _o_sv = 14'b10010101000110;
      11'b11000000110:
        _o_sv = 14'b10010101001100;
      11'b11000000111:
        _o_sv = 14'b10010101010010;
      11'b11000001000:
        _o_sv = 14'b10010101011000;
      11'b11000001001:
        _o_sv = 14'b10010101011110;
      11'b11000001010:
        _o_sv = 14'b10010101100100;
      11'b11000001011:
        _o_sv = 14'b10010101101010;
      11'b11000001100:
        _o_sv = 14'b10010101110000;
      11'b11000001101:
        _o_sv = 14'b10010101110110;
      11'b11000001110:
        _o_sv = 14'b10010101111100;
      11'b11000001111:
        _o_sv = 14'b10010110000010;
      11'b11000010000:
        _o_sv = 14'b10010110001000;
      11'b11000010001:
        _o_sv = 14'b10010110001110;
      11'b11000010010:
        _o_sv = 14'b10010110010100;
      11'b11000010011:
        _o_sv = 14'b10010110011010;
      11'b11000010100:
        _o_sv = 14'b10010110100000;
      11'b11000010101:
        _o_sv = 14'b10010110100110;
      11'b11000010110:
        _o_sv = 14'b10010110101100;
      11'b11000010111:
        _o_sv = 14'b10010110110010;
      11'b11000011000:
        _o_sv = 14'b10010110111000;
      11'b11000011001:
        _o_sv = 14'b10010110111110;
      11'b11000011010:
        _o_sv = 14'b10010111000100;
      11'b11000011011:
        _o_sv = 14'b10010111001010;
      11'b11000011100:
        _o_sv = 14'b10010111010000;
      11'b11000011101:
        _o_sv = 14'b10010111010110;
      11'b11000011110:
        _o_sv = 14'b10010111011100;
      11'b11000011111:
        _o_sv = 14'b10010111100010;
      11'b11000100000:
        _o_sv = 14'b10010111101000;
      11'b11000100001:
        _o_sv = 14'b10010111101110;
      11'b11000100010:
        _o_sv = 14'b10010111110100;
      11'b11000100011:
        _o_sv = 14'b10010111111010;
      11'b11000100100:
        _o_sv = 14'b10011000000000;
      11'b11000100101:
        _o_sv = 14'b10011000000110;
      11'b11000100110:
        _o_sv = 14'b10011000001100;
      11'b11000100111:
        _o_sv = 14'b10011000010010;
      11'b11000101000:
        _o_sv = 14'b10011000011000;
      11'b11000101001:
        _o_sv = 14'b10011000011110;
      11'b11000101010:
        _o_sv = 14'b10011000100100;
      11'b11000101011:
        _o_sv = 14'b10011000101010;
      11'b11000101100:
        _o_sv = 14'b10011000110000;
      11'b11000101101:
        _o_sv = 14'b10011000110110;
      11'b11000101110:
        _o_sv = 14'b10011000111100;
      11'b11000101111:
        _o_sv = 14'b10011001000010;
      11'b11000110000:
        _o_sv = 14'b10011001001000;
      11'b11000110001:
        _o_sv = 14'b10011001001110;
      11'b11000110010:
        _o_sv = 14'b10011001010100;
      11'b11000110011:
        _o_sv = 14'b10011001011010;
      11'b11000110100:
        _o_sv = 14'b10011001100000;
      11'b11000110101:
        _o_sv = 14'b10011001100110;
      11'b11000110110:
        _o_sv = 14'b10011001101100;
      11'b11000110111:
        _o_sv = 14'b10011001110010;
      11'b11000111000:
        _o_sv = 14'b10011001111000;
      11'b11000111001:
        _o_sv = 14'b10011001111110;
      11'b11000111010:
        _o_sv = 14'b10011010000100;
      11'b11000111011:
        _o_sv = 14'b10011010001010;
      11'b11000111100:
        _o_sv = 14'b10011010010000;
      11'b11000111101:
        _o_sv = 14'b10011010010110;
      11'b11000111110:
        _o_sv = 14'b10011010011100;
      11'b11000111111:
        _o_sv = 14'b10011010100010;
      11'b11001000000:
        _o_sv = 14'b10011010101000;
      11'b11001000001:
        _o_sv = 14'b10011010101110;
      11'b11001000010:
        _o_sv = 14'b10011010110100;
      11'b11001000011:
        _o_sv = 14'b10011010111010;
      11'b11001000100:
        _o_sv = 14'b10011011000000;
      11'b11001000101:
        _o_sv = 14'b10011011000110;
      11'b11001000110:
        _o_sv = 14'b10011011001100;
      11'b11001000111:
        _o_sv = 14'b10011011010010;
      11'b11001001000:
        _o_sv = 14'b10011011011000;
      11'b11001001001:
        _o_sv = 14'b10011011011110;
      11'b11001001010:
        _o_sv = 14'b10011011100100;
      11'b11001001011:
        _o_sv = 14'b10011011101001;
      11'b11001001100:
        _o_sv = 14'b10011011101111;
      11'b11001001101:
        _o_sv = 14'b10011011110101;
      11'b11001001110:
        _o_sv = 14'b10011011111011;
      11'b11001001111:
        _o_sv = 14'b10011100000001;
      11'b11001010000:
        _o_sv = 14'b10011100000111;
      11'b11001010001:
        _o_sv = 14'b10011100001101;
      11'b11001010010:
        _o_sv = 14'b10011100010011;
      11'b11001010011:
        _o_sv = 14'b10011100011001;
      11'b11001010100:
        _o_sv = 14'b10011100011111;
      11'b11001010101:
        _o_sv = 14'b10011100100101;
      11'b11001010110:
        _o_sv = 14'b10011100101011;
      11'b11001010111:
        _o_sv = 14'b10011100110001;
      11'b11001011000:
        _o_sv = 14'b10011100110111;
      11'b11001011001:
        _o_sv = 14'b10011100111101;
      11'b11001011010:
        _o_sv = 14'b10011101000011;
      11'b11001011011:
        _o_sv = 14'b10011101001001;
      11'b11001011100:
        _o_sv = 14'b10011101001111;
      11'b11001011101:
        _o_sv = 14'b10011101010101;
      11'b11001011110:
        _o_sv = 14'b10011101011011;
      11'b11001011111:
        _o_sv = 14'b10011101100001;
      11'b11001100000:
        _o_sv = 14'b10011101100111;
      11'b11001100001:
        _o_sv = 14'b10011101101101;
      11'b11001100010:
        _o_sv = 14'b10011101110011;
      11'b11001100011:
        _o_sv = 14'b10011101111001;
      11'b11001100100:
        _o_sv = 14'b10011101111111;
      11'b11001100101:
        _o_sv = 14'b10011110000101;
      11'b11001100110:
        _o_sv = 14'b10011110001011;
      11'b11001100111:
        _o_sv = 14'b10011110010001;
      11'b11001101000:
        _o_sv = 14'b10011110010111;
      11'b11001101001:
        _o_sv = 14'b10011110011101;
      11'b11001101010:
        _o_sv = 14'b10011110100011;
      11'b11001101011:
        _o_sv = 14'b10011110101001;
      11'b11001101100:
        _o_sv = 14'b10011110101111;
      11'b11001101101:
        _o_sv = 14'b10011110110101;
      11'b11001101110:
        _o_sv = 14'b10011110111011;
      11'b11001101111:
        _o_sv = 14'b10011111000001;
      11'b11001110000:
        _o_sv = 14'b10011111000111;
      11'b11001110001:
        _o_sv = 14'b10011111001101;
      11'b11001110010:
        _o_sv = 14'b10011111010011;
      11'b11001110011:
        _o_sv = 14'b10011111011001;
      11'b11001110100:
        _o_sv = 14'b10011111011111;
      11'b11001110101:
        _o_sv = 14'b10011111100101;
      11'b11001110110:
        _o_sv = 14'b10011111101011;
      11'b11001110111:
        _o_sv = 14'b10011111110001;
      11'b11001111000:
        _o_sv = 14'b10011111110110;
      11'b11001111001:
        _o_sv = 14'b10011111111100;
      11'b11001111010:
        _o_sv = 14'b10100000000010;
      11'b11001111011:
        _o_sv = 14'b10100000001000;
      11'b11001111100:
        _o_sv = 14'b10100000001110;
      11'b11001111101:
        _o_sv = 14'b10100000010100;
      11'b11001111110:
        _o_sv = 14'b10100000011010;
      11'b11001111111:
        _o_sv = 14'b10100000100000;
      11'b11010000000:
        _o_sv = 14'b10100000100110;
      11'b11010000001:
        _o_sv = 14'b10100000101100;
      11'b11010000010:
        _o_sv = 14'b10100000110010;
      11'b11010000011:
        _o_sv = 14'b10100000111000;
      11'b11010000100:
        _o_sv = 14'b10100000111110;
      11'b11010000101:
        _o_sv = 14'b10100001000100;
      11'b11010000110:
        _o_sv = 14'b10100001001010;
      11'b11010000111:
        _o_sv = 14'b10100001010000;
      11'b11010001000:
        _o_sv = 14'b10100001010110;
      11'b11010001001:
        _o_sv = 14'b10100001011100;
      11'b11010001010:
        _o_sv = 14'b10100001100010;
      11'b11010001011:
        _o_sv = 14'b10100001101000;
      11'b11010001100:
        _o_sv = 14'b10100001101110;
      11'b11010001101:
        _o_sv = 14'b10100001110100;
      11'b11010001110:
        _o_sv = 14'b10100001111010;
      11'b11010001111:
        _o_sv = 14'b10100010000000;
      11'b11010010000:
        _o_sv = 14'b10100010000110;
      11'b11010010001:
        _o_sv = 14'b10100010001100;
      11'b11010010010:
        _o_sv = 14'b10100010010010;
      11'b11010010011:
        _o_sv = 14'b10100010011000;
      11'b11010010100:
        _o_sv = 14'b10100010011101;
      11'b11010010101:
        _o_sv = 14'b10100010100011;
      11'b11010010110:
        _o_sv = 14'b10100010101001;
      11'b11010010111:
        _o_sv = 14'b10100010101111;
      11'b11010011000:
        _o_sv = 14'b10100010110101;
      11'b11010011001:
        _o_sv = 14'b10100010111011;
      11'b11010011010:
        _o_sv = 14'b10100011000001;
      11'b11010011011:
        _o_sv = 14'b10100011000111;
      11'b11010011100:
        _o_sv = 14'b10100011001101;
      11'b11010011101:
        _o_sv = 14'b10100011010011;
      11'b11010011110:
        _o_sv = 14'b10100011011001;
      11'b11010011111:
        _o_sv = 14'b10100011011111;
      11'b11010100000:
        _o_sv = 14'b10100011100101;
      11'b11010100001:
        _o_sv = 14'b10100011101011;
      11'b11010100010:
        _o_sv = 14'b10100011110001;
      11'b11010100011:
        _o_sv = 14'b10100011110111;
      11'b11010100100:
        _o_sv = 14'b10100011111101;
      11'b11010100101:
        _o_sv = 14'b10100100000011;
      11'b11010100110:
        _o_sv = 14'b10100100001001;
      11'b11010100111:
        _o_sv = 14'b10100100001111;
      11'b11010101000:
        _o_sv = 14'b10100100010101;
      11'b11010101001:
        _o_sv = 14'b10100100011011;
      11'b11010101010:
        _o_sv = 14'b10100100100000;
      11'b11010101011:
        _o_sv = 14'b10100100100110;
      11'b11010101100:
        _o_sv = 14'b10100100101100;
      11'b11010101101:
        _o_sv = 14'b10100100110010;
      11'b11010101110:
        _o_sv = 14'b10100100111000;
      11'b11010101111:
        _o_sv = 14'b10100100111110;
      11'b11010110000:
        _o_sv = 14'b10100101000100;
      11'b11010110001:
        _o_sv = 14'b10100101001010;
      11'b11010110010:
        _o_sv = 14'b10100101010000;
      11'b11010110011:
        _o_sv = 14'b10100101010110;
      11'b11010110100:
        _o_sv = 14'b10100101011100;
      11'b11010110101:
        _o_sv = 14'b10100101100010;
      11'b11010110110:
        _o_sv = 14'b10100101101000;
      11'b11010110111:
        _o_sv = 14'b10100101101110;
      11'b11010111000:
        _o_sv = 14'b10100101110100;
      11'b11010111001:
        _o_sv = 14'b10100101111010;
      11'b11010111010:
        _o_sv = 14'b10100110000000;
      11'b11010111011:
        _o_sv = 14'b10100110000110;
      11'b11010111100:
        _o_sv = 14'b10100110001011;
      11'b11010111101:
        _o_sv = 14'b10100110010001;
      11'b11010111110:
        _o_sv = 14'b10100110010111;
      11'b11010111111:
        _o_sv = 14'b10100110011101;
      11'b11011000000:
        _o_sv = 14'b10100110100011;
      11'b11011000001:
        _o_sv = 14'b10100110101001;
      11'b11011000010:
        _o_sv = 14'b10100110101111;
      11'b11011000011:
        _o_sv = 14'b10100110110101;
      11'b11011000100:
        _o_sv = 14'b10100110111011;
      11'b11011000101:
        _o_sv = 14'b10100111000001;
      11'b11011000110:
        _o_sv = 14'b10100111000111;
      11'b11011000111:
        _o_sv = 14'b10100111001101;
      11'b11011001000:
        _o_sv = 14'b10100111010011;
      11'b11011001001:
        _o_sv = 14'b10100111011001;
      11'b11011001010:
        _o_sv = 14'b10100111011111;
      11'b11011001011:
        _o_sv = 14'b10100111100101;
      11'b11011001100:
        _o_sv = 14'b10100111101011;
      11'b11011001101:
        _o_sv = 14'b10100111110000;
      11'b11011001110:
        _o_sv = 14'b10100111110110;
      11'b11011001111:
        _o_sv = 14'b10100111111100;
      11'b11011010000:
        _o_sv = 14'b10101000000010;
      11'b11011010001:
        _o_sv = 14'b10101000001000;
      11'b11011010010:
        _o_sv = 14'b10101000001110;
      11'b11011010011:
        _o_sv = 14'b10101000010100;
      11'b11011010100:
        _o_sv = 14'b10101000011010;
      11'b11011010101:
        _o_sv = 14'b10101000100000;
      11'b11011010110:
        _o_sv = 14'b10101000100110;
      11'b11011010111:
        _o_sv = 14'b10101000101100;
      11'b11011011000:
        _o_sv = 14'b10101000110010;
      11'b11011011001:
        _o_sv = 14'b10101000111000;
      11'b11011011010:
        _o_sv = 14'b10101000111110;
      11'b11011011011:
        _o_sv = 14'b10101001000100;
      11'b11011011100:
        _o_sv = 14'b10101001001001;
      11'b11011011101:
        _o_sv = 14'b10101001001111;
      11'b11011011110:
        _o_sv = 14'b10101001010101;
      11'b11011011111:
        _o_sv = 14'b10101001011011;
      11'b11011100000:
        _o_sv = 14'b10101001100001;
      11'b11011100001:
        _o_sv = 14'b10101001100111;
      11'b11011100010:
        _o_sv = 14'b10101001101101;
      11'b11011100011:
        _o_sv = 14'b10101001110011;
      11'b11011100100:
        _o_sv = 14'b10101001111001;
      11'b11011100101:
        _o_sv = 14'b10101001111111;
      11'b11011100110:
        _o_sv = 14'b10101010000101;
      11'b11011100111:
        _o_sv = 14'b10101010001011;
      11'b11011101000:
        _o_sv = 14'b10101010010001;
      11'b11011101001:
        _o_sv = 14'b10101010010111;
      11'b11011101010:
        _o_sv = 14'b10101010011100;
      11'b11011101011:
        _o_sv = 14'b10101010100010;
      11'b11011101100:
        _o_sv = 14'b10101010101000;
      11'b11011101101:
        _o_sv = 14'b10101010101110;
      11'b11011101110:
        _o_sv = 14'b10101010110100;
      11'b11011101111:
        _o_sv = 14'b10101010111010;
      11'b11011110000:
        _o_sv = 14'b10101011000000;
      11'b11011110001:
        _o_sv = 14'b10101011000110;
      11'b11011110010:
        _o_sv = 14'b10101011001100;
      11'b11011110011:
        _o_sv = 14'b10101011010010;
      11'b11011110100:
        _o_sv = 14'b10101011011000;
      11'b11011110101:
        _o_sv = 14'b10101011011110;
      11'b11011110110:
        _o_sv = 14'b10101011100100;
      11'b11011110111:
        _o_sv = 14'b10101011101001;
      11'b11011111000:
        _o_sv = 14'b10101011101111;
      11'b11011111001:
        _o_sv = 14'b10101011110101;
      11'b11011111010:
        _o_sv = 14'b10101011111011;
      11'b11011111011:
        _o_sv = 14'b10101100000001;
      11'b11011111100:
        _o_sv = 14'b10101100000111;
      11'b11011111101:
        _o_sv = 14'b10101100001101;
      11'b11011111110:
        _o_sv = 14'b10101100010011;
      11'b11011111111:
        _o_sv = 14'b10101100011001;
      11'b11100000000:
        _o_sv = 14'b10101100011111;
      11'b11100000001:
        _o_sv = 14'b10101100100101;
      11'b11100000010:
        _o_sv = 14'b10101100101011;
      11'b11100000011:
        _o_sv = 14'b10101100110000;
      11'b11100000100:
        _o_sv = 14'b10101100110110;
      11'b11100000101:
        _o_sv = 14'b10101100111100;
      11'b11100000110:
        _o_sv = 14'b10101101000010;
      11'b11100000111:
        _o_sv = 14'b10101101001000;
      11'b11100001000:
        _o_sv = 14'b10101101001110;
      11'b11100001001:
        _o_sv = 14'b10101101010100;
      11'b11100001010:
        _o_sv = 14'b10101101011010;
      11'b11100001011:
        _o_sv = 14'b10101101100000;
      11'b11100001100:
        _o_sv = 14'b10101101100110;
      11'b11100001101:
        _o_sv = 14'b10101101101100;
      11'b11100001110:
        _o_sv = 14'b10101101110001;
      11'b11100001111:
        _o_sv = 14'b10101101110111;
      11'b11100010000:
        _o_sv = 14'b10101101111101;
      11'b11100010001:
        _o_sv = 14'b10101110000011;
      11'b11100010010:
        _o_sv = 14'b10101110001001;
      11'b11100010011:
        _o_sv = 14'b10101110001111;
      11'b11100010100:
        _o_sv = 14'b10101110010101;
      11'b11100010101:
        _o_sv = 14'b10101110011011;
      11'b11100010110:
        _o_sv = 14'b10101110100001;
      11'b11100010111:
        _o_sv = 14'b10101110100111;
      11'b11100011000:
        _o_sv = 14'b10101110101101;
      11'b11100011001:
        _o_sv = 14'b10101110110010;
      11'b11100011010:
        _o_sv = 14'b10101110111000;
      11'b11100011011:
        _o_sv = 14'b10101110111110;
      11'b11100011100:
        _o_sv = 14'b10101111000100;
      11'b11100011101:
        _o_sv = 14'b10101111001010;
      11'b11100011110:
        _o_sv = 14'b10101111010000;
      11'b11100011111:
        _o_sv = 14'b10101111010110;
      11'b11100100000:
        _o_sv = 14'b10101111011100;
      11'b11100100001:
        _o_sv = 14'b10101111100010;
      11'b11100100010:
        _o_sv = 14'b10101111101000;
      11'b11100100011:
        _o_sv = 14'b10101111101110;
      11'b11100100100:
        _o_sv = 14'b10101111110011;
      11'b11100100101:
        _o_sv = 14'b10101111111001;
      11'b11100100110:
        _o_sv = 14'b10101111111111;
      11'b11100100111:
        _o_sv = 14'b10110000000101;
      11'b11100101000:
        _o_sv = 14'b10110000001011;
      11'b11100101001:
        _o_sv = 14'b10110000010001;
      11'b11100101010:
        _o_sv = 14'b10110000010111;
      11'b11100101011:
        _o_sv = 14'b10110000011101;
      11'b11100101100:
        _o_sv = 14'b10110000100011;
      11'b11100101101:
        _o_sv = 14'b10110000101001;
      11'b11100101110:
        _o_sv = 14'b10110000101110;
      11'b11100101111:
        _o_sv = 14'b10110000110100;
      11'b11100110000:
        _o_sv = 14'b10110000111010;
      11'b11100110001:
        _o_sv = 14'b10110001000000;
      11'b11100110010:
        _o_sv = 14'b10110001000110;
      11'b11100110011:
        _o_sv = 14'b10110001001100;
      11'b11100110100:
        _o_sv = 14'b10110001010010;
      11'b11100110101:
        _o_sv = 14'b10110001011000;
      11'b11100110110:
        _o_sv = 14'b10110001011110;
      11'b11100110111:
        _o_sv = 14'b10110001100011;
      11'b11100111000:
        _o_sv = 14'b10110001101001;
      11'b11100111001:
        _o_sv = 14'b10110001101111;
      11'b11100111010:
        _o_sv = 14'b10110001110101;
      11'b11100111011:
        _o_sv = 14'b10110001111011;
      11'b11100111100:
        _o_sv = 14'b10110010000001;
      11'b11100111101:
        _o_sv = 14'b10110010000111;
      11'b11100111110:
        _o_sv = 14'b10110010001101;
      11'b11100111111:
        _o_sv = 14'b10110010010011;
      11'b11101000000:
        _o_sv = 14'b10110010011000;
      11'b11101000001:
        _o_sv = 14'b10110010011110;
      11'b11101000010:
        _o_sv = 14'b10110010100100;
      11'b11101000011:
        _o_sv = 14'b10110010101010;
      11'b11101000100:
        _o_sv = 14'b10110010110000;
      11'b11101000101:
        _o_sv = 14'b10110010110110;
      11'b11101000110:
        _o_sv = 14'b10110010111100;
      11'b11101000111:
        _o_sv = 14'b10110011000010;
      11'b11101001000:
        _o_sv = 14'b10110011001000;
      11'b11101001001:
        _o_sv = 14'b10110011001101;
      11'b11101001010:
        _o_sv = 14'b10110011010011;
      11'b11101001011:
        _o_sv = 14'b10110011011001;
      11'b11101001100:
        _o_sv = 14'b10110011011111;
      11'b11101001101:
        _o_sv = 14'b10110011100101;
      11'b11101001110:
        _o_sv = 14'b10110011101011;
      11'b11101001111:
        _o_sv = 14'b10110011110001;
      11'b11101010000:
        _o_sv = 14'b10110011110111;
      11'b11101010001:
        _o_sv = 14'b10110011111101;
      11'b11101010010:
        _o_sv = 14'b10110100000010;
      11'b11101010011:
        _o_sv = 14'b10110100001000;
      11'b11101010100:
        _o_sv = 14'b10110100001110;
      11'b11101010101:
        _o_sv = 14'b10110100010100;
      11'b11101010110:
        _o_sv = 14'b10110100011010;
      11'b11101010111:
        _o_sv = 14'b10110100100000;
      11'b11101011000:
        _o_sv = 14'b10110100100110;
      11'b11101011001:
        _o_sv = 14'b10110100101100;
      11'b11101011010:
        _o_sv = 14'b10110100110001;
      11'b11101011011:
        _o_sv = 14'b10110100110111;
      11'b11101011100:
        _o_sv = 14'b10110100111101;
      11'b11101011101:
        _o_sv = 14'b10110101000011;
      11'b11101011110:
        _o_sv = 14'b10110101001001;
      11'b11101011111:
        _o_sv = 14'b10110101001111;
      11'b11101100000:
        _o_sv = 14'b10110101010101;
      11'b11101100001:
        _o_sv = 14'b10110101011011;
      11'b11101100010:
        _o_sv = 14'b10110101100000;
      11'b11101100011:
        _o_sv = 14'b10110101100110;
      11'b11101100100:
        _o_sv = 14'b10110101101100;
      11'b11101100101:
        _o_sv = 14'b10110101110010;
      11'b11101100110:
        _o_sv = 14'b10110101111000;
      11'b11101100111:
        _o_sv = 14'b10110101111110;
      11'b11101101000:
        _o_sv = 14'b10110110000100;
      11'b11101101001:
        _o_sv = 14'b10110110001010;
      11'b11101101010:
        _o_sv = 14'b10110110001111;
      11'b11101101011:
        _o_sv = 14'b10110110010101;
      11'b11101101100:
        _o_sv = 14'b10110110011011;
      11'b11101101101:
        _o_sv = 14'b10110110100001;
      11'b11101101110:
        _o_sv = 14'b10110110100111;
      11'b11101101111:
        _o_sv = 14'b10110110101101;
      11'b11101110000:
        _o_sv = 14'b10110110110011;
      11'b11101110001:
        _o_sv = 14'b10110110111001;
      11'b11101110010:
        _o_sv = 14'b10110110111110;
      11'b11101110011:
        _o_sv = 14'b10110111000100;
      11'b11101110100:
        _o_sv = 14'b10110111001010;
      11'b11101110101:
        _o_sv = 14'b10110111010000;
      11'b11101110110:
        _o_sv = 14'b10110111010110;
      11'b11101110111:
        _o_sv = 14'b10110111011100;
      11'b11101111000:
        _o_sv = 14'b10110111100010;
      11'b11101111001:
        _o_sv = 14'b10110111100111;
      11'b11101111010:
        _o_sv = 14'b10110111101101;
      11'b11101111011:
        _o_sv = 14'b10110111110011;
      11'b11101111100:
        _o_sv = 14'b10110111111001;
      11'b11101111101:
        _o_sv = 14'b10110111111111;
      11'b11101111110:
        _o_sv = 14'b10111000000101;
      11'b11101111111:
        _o_sv = 14'b10111000001011;
      11'b11110000000:
        _o_sv = 14'b10111000010001;
      11'b11110000001:
        _o_sv = 14'b10111000010110;
      11'b11110000010:
        _o_sv = 14'b10111000011100;
      11'b11110000011:
        _o_sv = 14'b10111000100010;
      11'b11110000100:
        _o_sv = 14'b10111000101000;
      11'b11110000101:
        _o_sv = 14'b10111000101110;
      11'b11110000110:
        _o_sv = 14'b10111000110100;
      11'b11110000111:
        _o_sv = 14'b10111000111010;
      11'b11110001000:
        _o_sv = 14'b10111000111111;
      11'b11110001001:
        _o_sv = 14'b10111001000101;
      11'b11110001010:
        _o_sv = 14'b10111001001011;
      11'b11110001011:
        _o_sv = 14'b10111001010001;
      11'b11110001100:
        _o_sv = 14'b10111001010111;
      11'b11110001101:
        _o_sv = 14'b10111001011101;
      11'b11110001110:
        _o_sv = 14'b10111001100011;
      11'b11110001111:
        _o_sv = 14'b10111001101000;
      11'b11110010000:
        _o_sv = 14'b10111001101110;
      11'b11110010001:
        _o_sv = 14'b10111001110100;
      11'b11110010010:
        _o_sv = 14'b10111001111010;
      11'b11110010011:
        _o_sv = 14'b10111010000000;
      11'b11110010100:
        _o_sv = 14'b10111010000110;
      11'b11110010101:
        _o_sv = 14'b10111010001100;
      11'b11110010110:
        _o_sv = 14'b10111010010001;
      11'b11110010111:
        _o_sv = 14'b10111010010111;
      11'b11110011000:
        _o_sv = 14'b10111010011101;
      11'b11110011001:
        _o_sv = 14'b10111010100011;
      11'b11110011010:
        _o_sv = 14'b10111010101001;
      11'b11110011011:
        _o_sv = 14'b10111010101111;
      11'b11110011100:
        _o_sv = 14'b10111010110101;
      11'b11110011101:
        _o_sv = 14'b10111010111010;
      11'b11110011110:
        _o_sv = 14'b10111011000000;
      11'b11110011111:
        _o_sv = 14'b10111011000110;
      11'b11110100000:
        _o_sv = 14'b10111011001100;
      11'b11110100001:
        _o_sv = 14'b10111011010010;
      11'b11110100010:
        _o_sv = 14'b10111011011000;
      11'b11110100011:
        _o_sv = 14'b10111011011101;
      11'b11110100100:
        _o_sv = 14'b10111011100011;
      11'b11110100101:
        _o_sv = 14'b10111011101001;
      11'b11110100110:
        _o_sv = 14'b10111011101111;
      11'b11110100111:
        _o_sv = 14'b10111011110101;
      11'b11110101000:
        _o_sv = 14'b10111011111011;
      11'b11110101001:
        _o_sv = 14'b10111100000001;
      11'b11110101010:
        _o_sv = 14'b10111100000110;
      11'b11110101011:
        _o_sv = 14'b10111100001100;
      11'b11110101100:
        _o_sv = 14'b10111100010010;
      11'b11110101101:
        _o_sv = 14'b10111100011000;
      11'b11110101110:
        _o_sv = 14'b10111100011110;
      11'b11110101111:
        _o_sv = 14'b10111100100100;
      11'b11110110000:
        _o_sv = 14'b10111100101001;
      11'b11110110001:
        _o_sv = 14'b10111100101111;
      11'b11110110010:
        _o_sv = 14'b10111100110101;
      11'b11110110011:
        _o_sv = 14'b10111100111011;
      11'b11110110100:
        _o_sv = 14'b10111101000001;
      11'b11110110101:
        _o_sv = 14'b10111101000111;
      11'b11110110110:
        _o_sv = 14'b10111101001100;
      11'b11110110111:
        _o_sv = 14'b10111101010010;
      11'b11110111000:
        _o_sv = 14'b10111101011000;
      11'b11110111001:
        _o_sv = 14'b10111101011110;
      11'b11110111010:
        _o_sv = 14'b10111101100100;
      11'b11110111011:
        _o_sv = 14'b10111101101010;
      11'b11110111100:
        _o_sv = 14'b10111101101111;
      11'b11110111101:
        _o_sv = 14'b10111101110101;
      11'b11110111110:
        _o_sv = 14'b10111101111011;
      11'b11110111111:
        _o_sv = 14'b10111110000001;
      11'b11111000000:
        _o_sv = 14'b10111110000111;
      11'b11111000001:
        _o_sv = 14'b10111110001101;
      11'b11111000010:
        _o_sv = 14'b10111110010010;
      11'b11111000011:
        _o_sv = 14'b10111110011000;
      11'b11111000100:
        _o_sv = 14'b10111110011110;
      11'b11111000101:
        _o_sv = 14'b10111110100100;
      11'b11111000110:
        _o_sv = 14'b10111110101010;
      11'b11111000111:
        _o_sv = 14'b10111110110000;
      11'b11111001000:
        _o_sv = 14'b10111110110101;
      11'b11111001001:
        _o_sv = 14'b10111110111011;
      11'b11111001010:
        _o_sv = 14'b10111111000001;
      11'b11111001011:
        _o_sv = 14'b10111111000111;
      11'b11111001100:
        _o_sv = 14'b10111111001101;
      11'b11111001101:
        _o_sv = 14'b10111111010011;
      11'b11111001110:
        _o_sv = 14'b10111111011000;
      11'b11111001111:
        _o_sv = 14'b10111111011110;
      11'b11111010000:
        _o_sv = 14'b10111111100100;
      11'b11111010001:
        _o_sv = 14'b10111111101010;
      11'b11111010010:
        _o_sv = 14'b10111111110000;
      11'b11111010011:
        _o_sv = 14'b10111111110110;
      11'b11111010100:
        _o_sv = 14'b10111111111011;
      11'b11111010101:
        _o_sv = 14'b11000000000001;
      11'b11111010110:
        _o_sv = 14'b11000000000111;
      11'b11111010111:
        _o_sv = 14'b11000000001101;
      11'b11111011000:
        _o_sv = 14'b11000000010011;
      11'b11111011001:
        _o_sv = 14'b11000000011001;
      11'b11111011010:
        _o_sv = 14'b11000000011110;
      11'b11111011011:
        _o_sv = 14'b11000000100100;
      11'b11111011100:
        _o_sv = 14'b11000000101010;
      11'b11111011101:
        _o_sv = 14'b11000000110000;
      11'b11111011110:
        _o_sv = 14'b11000000110110;
      11'b11111011111:
        _o_sv = 14'b11000000111011;
      11'b11111100000:
        _o_sv = 14'b11000001000001;
      11'b11111100001:
        _o_sv = 14'b11000001000111;
      11'b11111100010:
        _o_sv = 14'b11000001001101;
      11'b11111100011:
        _o_sv = 14'b11000001010011;
      11'b11111100100:
        _o_sv = 14'b11000001011001;
      11'b11111100101:
        _o_sv = 14'b11000001011110;
      11'b11111100110:
        _o_sv = 14'b11000001100100;
      11'b11111100111:
        _o_sv = 14'b11000001101010;
      11'b11111101000:
        _o_sv = 14'b11000001110000;
      11'b11111101001:
        _o_sv = 14'b11000001110110;
      11'b11111101010:
        _o_sv = 14'b11000001111011;
      11'b11111101011:
        _o_sv = 14'b11000010000001;
      11'b11111101100:
        _o_sv = 14'b11000010000111;
      11'b11111101101:
        _o_sv = 14'b11000010001101;
      11'b11111101110:
        _o_sv = 14'b11000010010011;
      11'b11111101111:
        _o_sv = 14'b11000010011001;
      11'b11111110000:
        _o_sv = 14'b11000010011110;
      11'b11111110001:
        _o_sv = 14'b11000010100100;
      11'b11111110010:
        _o_sv = 14'b11000010101010;
      11'b11111110011:
        _o_sv = 14'b11000010110000;
      11'b11111110100:
        _o_sv = 14'b11000010110110;
      11'b11111110101:
        _o_sv = 14'b11000010111011;
      11'b11111110110:
        _o_sv = 14'b11000011000001;
      11'b11111110111:
        _o_sv = 14'b11000011000111;
      11'b11111111000:
        _o_sv = 14'b11000011001101;
      11'b11111111001:
        _o_sv = 14'b11000011010011;
      11'b11111111010:
        _o_sv = 14'b11000011011000;
      11'b11111111011:
        _o_sv = 14'b11000011011110;
      11'b11111111100:
        _o_sv = 14'b11000011100100;
      11'b11111111101:
        _o_sv = 14'b11000011101010;
      11'b11111111110:
        _o_sv = 14'b11000011110000;
      11'b11111111111:
        _o_sv = 14'b11000011110101;
      12'b100000000000:
        _o_sv = 14'b11000011111011;
      12'b100000000001:
        _o_sv = 14'b11000100000001;
      12'b100000000010:
        _o_sv = 14'b11000100000111;
      12'b100000000011:
        _o_sv = 14'b11000100001101;
      12'b100000000100:
        _o_sv = 14'b11000100010010;
      12'b100000000101:
        _o_sv = 14'b11000100011000;
      12'b100000000110:
        _o_sv = 14'b11000100011110;
      12'b100000000111:
        _o_sv = 14'b11000100100100;
      12'b100000001000:
        _o_sv = 14'b11000100101010;
      12'b100000001001:
        _o_sv = 14'b11000100101111;
      12'b100000001010:
        _o_sv = 14'b11000100110101;
      12'b100000001011:
        _o_sv = 14'b11000100111011;
      12'b100000001100:
        _o_sv = 14'b11000101000001;
      12'b100000001101:
        _o_sv = 14'b11000101000111;
      12'b100000001110:
        _o_sv = 14'b11000101001100;
      12'b100000001111:
        _o_sv = 14'b11000101010010;
      12'b100000010000:
        _o_sv = 14'b11000101011000;
      12'b100000010001:
        _o_sv = 14'b11000101011110;
      12'b100000010010:
        _o_sv = 14'b11000101100100;
      12'b100000010011:
        _o_sv = 14'b11000101101001;
      12'b100000010100:
        _o_sv = 14'b11000101101111;
      12'b100000010101:
        _o_sv = 14'b11000101110101;
      12'b100000010110:
        _o_sv = 14'b11000101111011;
      12'b100000010111:
        _o_sv = 14'b11000110000001;
      12'b100000011000:
        _o_sv = 14'b11000110000110;
      12'b100000011001:
        _o_sv = 14'b11000110001100;
      12'b100000011010:
        _o_sv = 14'b11000110010010;
      12'b100000011011:
        _o_sv = 14'b11000110011000;
      12'b100000011100:
        _o_sv = 14'b11000110011110;
      12'b100000011101:
        _o_sv = 14'b11000110100011;
      12'b100000011110:
        _o_sv = 14'b11000110101001;
      12'b100000011111:
        _o_sv = 14'b11000110101111;
      12'b100000100000:
        _o_sv = 14'b11000110110101;
      12'b100000100001:
        _o_sv = 14'b11000110111011;
      12'b100000100010:
        _o_sv = 14'b11000111000000;
      12'b100000100011:
        _o_sv = 14'b11000111000110;
      12'b100000100100:
        _o_sv = 14'b11000111001100;
      12'b100000100101:
        _o_sv = 14'b11000111010010;
      12'b100000100110:
        _o_sv = 14'b11000111011000;
      12'b100000100111:
        _o_sv = 14'b11000111011101;
      12'b100000101000:
        _o_sv = 14'b11000111100011;
      12'b100000101001:
        _o_sv = 14'b11000111101001;
      12'b100000101010:
        _o_sv = 14'b11000111101111;
      12'b100000101011:
        _o_sv = 14'b11000111110100;
      12'b100000101100:
        _o_sv = 14'b11000111111010;
      12'b100000101101:
        _o_sv = 14'b11001000000000;
      12'b100000101110:
        _o_sv = 14'b11001000000110;
      12'b100000101111:
        _o_sv = 14'b11001000001100;
      12'b100000110000:
        _o_sv = 14'b11001000010001;
      12'b100000110001:
        _o_sv = 14'b11001000010111;
      12'b100000110010:
        _o_sv = 14'b11001000011101;
      12'b100000110011:
        _o_sv = 14'b11001000100011;
      12'b100000110100:
        _o_sv = 14'b11001000101000;
      12'b100000110101:
        _o_sv = 14'b11001000101110;
      12'b100000110110:
        _o_sv = 14'b11001000110100;
      12'b100000110111:
        _o_sv = 14'b11001000111010;
      12'b100000111000:
        _o_sv = 14'b11001001000000;
      12'b100000111001:
        _o_sv = 14'b11001001000101;
      12'b100000111010:
        _o_sv = 14'b11001001001011;
      12'b100000111011:
        _o_sv = 14'b11001001010001;
      12'b100000111100:
        _o_sv = 14'b11001001010111;
      12'b100000111101:
        _o_sv = 14'b11001001011101;
      12'b100000111110:
        _o_sv = 14'b11001001100010;
      12'b100000111111:
        _o_sv = 14'b11001001101000;
      12'b100001000000:
        _o_sv = 14'b11001001101110;
      12'b100001000001:
        _o_sv = 14'b11001001110100;
      12'b100001000010:
        _o_sv = 14'b11001001111001;
      12'b100001000011:
        _o_sv = 14'b11001001111111;
      12'b100001000100:
        _o_sv = 14'b11001010000101;
      12'b100001000101:
        _o_sv = 14'b11001010001011;
      12'b100001000110:
        _o_sv = 14'b11001010010000;
      12'b100001000111:
        _o_sv = 14'b11001010010110;
      12'b100001001000:
        _o_sv = 14'b11001010011100;
      12'b100001001001:
        _o_sv = 14'b11001010100010;
      12'b100001001010:
        _o_sv = 14'b11001010101000;
      12'b100001001011:
        _o_sv = 14'b11001010101101;
      12'b100001001100:
        _o_sv = 14'b11001010110011;
      12'b100001001101:
        _o_sv = 14'b11001010111001;
      12'b100001001110:
        _o_sv = 14'b11001010111111;
      12'b100001001111:
        _o_sv = 14'b11001011000100;
      12'b100001010000:
        _o_sv = 14'b11001011001010;
      12'b100001010001:
        _o_sv = 14'b11001011010000;
      12'b100001010010:
        _o_sv = 14'b11001011010110;
      12'b100001010011:
        _o_sv = 14'b11001011011011;
      12'b100001010100:
        _o_sv = 14'b11001011100001;
      12'b100001010101:
        _o_sv = 14'b11001011100111;
      12'b100001010110:
        _o_sv = 14'b11001011101101;
      12'b100001010111:
        _o_sv = 14'b11001011110011;
      12'b100001011000:
        _o_sv = 14'b11001011111000;
      12'b100001011001:
        _o_sv = 14'b11001011111110;
      12'b100001011010:
        _o_sv = 14'b11001100000100;
      12'b100001011011:
        _o_sv = 14'b11001100001010;
      12'b100001011100:
        _o_sv = 14'b11001100001111;
      12'b100001011101:
        _o_sv = 14'b11001100010101;
      12'b100001011110:
        _o_sv = 14'b11001100011011;
      12'b100001011111:
        _o_sv = 14'b11001100100001;
      12'b100001100000:
        _o_sv = 14'b11001100100110;
      12'b100001100001:
        _o_sv = 14'b11001100101100;
      12'b100001100010:
        _o_sv = 14'b11001100110010;
      12'b100001100011:
        _o_sv = 14'b11001100111000;
      12'b100001100100:
        _o_sv = 14'b11001100111101;
      12'b100001100101:
        _o_sv = 14'b11001101000011;
      12'b100001100110:
        _o_sv = 14'b11001101001001;
      12'b100001100111:
        _o_sv = 14'b11001101001111;
      12'b100001101000:
        _o_sv = 14'b11001101010100;
      12'b100001101001:
        _o_sv = 14'b11001101011010;
      12'b100001101010:
        _o_sv = 14'b11001101100000;
      12'b100001101011:
        _o_sv = 14'b11001101100110;
      12'b100001101100:
        _o_sv = 14'b11001101101011;
      12'b100001101101:
        _o_sv = 14'b11001101110001;
      12'b100001101110:
        _o_sv = 14'b11001101110111;
      12'b100001101111:
        _o_sv = 14'b11001101111101;
      12'b100001110000:
        _o_sv = 14'b11001110000010;
      12'b100001110001:
        _o_sv = 14'b11001110001000;
      12'b100001110010:
        _o_sv = 14'b11001110001110;
      12'b100001110011:
        _o_sv = 14'b11001110010100;
      12'b100001110100:
        _o_sv = 14'b11001110011001;
      12'b100001110101:
        _o_sv = 14'b11001110011111;
      12'b100001110110:
        _o_sv = 14'b11001110100101;
      12'b100001110111:
        _o_sv = 14'b11001110101011;
      12'b100001111000:
        _o_sv = 14'b11001110110000;
      12'b100001111001:
        _o_sv = 14'b11001110110110;
      12'b100001111010:
        _o_sv = 14'b11001110111100;
      12'b100001111011:
        _o_sv = 14'b11001111000010;
      12'b100001111100:
        _o_sv = 14'b11001111000111;
      12'b100001111101:
        _o_sv = 14'b11001111001101;
      12'b100001111110:
        _o_sv = 14'b11001111010011;
      12'b100001111111:
        _o_sv = 14'b11001111011001;
      12'b100010000000:
        _o_sv = 14'b11001111011110;
      12'b100010000001:
        _o_sv = 14'b11001111100100;
      12'b100010000010:
        _o_sv = 14'b11001111101010;
      12'b100010000011:
        _o_sv = 14'b11001111110000;
      12'b100010000100:
        _o_sv = 14'b11001111110101;
      12'b100010000101:
        _o_sv = 14'b11001111111011;
      12'b100010000110:
        _o_sv = 14'b11010000000001;
      12'b100010000111:
        _o_sv = 14'b11010000000111;
      12'b100010001000:
        _o_sv = 14'b11010000001100;
      12'b100010001001:
        _o_sv = 14'b11010000010010;
      12'b100010001010:
        _o_sv = 14'b11010000011000;
      12'b100010001011:
        _o_sv = 14'b11010000011110;
      12'b100010001100:
        _o_sv = 14'b11010000100011;
      12'b100010001101:
        _o_sv = 14'b11010000101001;
      12'b100010001110:
        _o_sv = 14'b11010000101111;
      12'b100010001111:
        _o_sv = 14'b11010000110101;
      12'b100010010000:
        _o_sv = 14'b11010000111010;
      12'b100010010001:
        _o_sv = 14'b11010001000000;
      12'b100010010010:
        _o_sv = 14'b11010001000110;
      12'b100010010011:
        _o_sv = 14'b11010001001011;
      12'b100010010100:
        _o_sv = 14'b11010001010001;
      12'b100010010101:
        _o_sv = 14'b11010001010111;
      12'b100010010110:
        _o_sv = 14'b11010001011101;
      12'b100010010111:
        _o_sv = 14'b11010001100010;
      12'b100010011000:
        _o_sv = 14'b11010001101000;
      12'b100010011001:
        _o_sv = 14'b11010001101110;
      12'b100010011010:
        _o_sv = 14'b11010001110100;
      12'b100010011011:
        _o_sv = 14'b11010001111001;
      12'b100010011100:
        _o_sv = 14'b11010001111111;
      12'b100010011101:
        _o_sv = 14'b11010010000101;
      12'b100010011110:
        _o_sv = 14'b11010010001011;
      12'b100010011111:
        _o_sv = 14'b11010010010000;
      12'b100010100000:
        _o_sv = 14'b11010010010110;
      12'b100010100001:
        _o_sv = 14'b11010010011100;
      12'b100010100010:
        _o_sv = 14'b11010010100001;
      12'b100010100011:
        _o_sv = 14'b11010010100111;
      12'b100010100100:
        _o_sv = 14'b11010010101101;
      12'b100010100101:
        _o_sv = 14'b11010010110011;
      12'b100010100110:
        _o_sv = 14'b11010010111000;
      12'b100010100111:
        _o_sv = 14'b11010010111110;
      12'b100010101000:
        _o_sv = 14'b11010011000100;
      12'b100010101001:
        _o_sv = 14'b11010011001010;
      12'b100010101010:
        _o_sv = 14'b11010011001111;
      12'b100010101011:
        _o_sv = 14'b11010011010101;
      12'b100010101100:
        _o_sv = 14'b11010011011011;
      12'b100010101101:
        _o_sv = 14'b11010011100000;
      12'b100010101110:
        _o_sv = 14'b11010011100110;
      12'b100010101111:
        _o_sv = 14'b11010011101100;
      12'b100010110000:
        _o_sv = 14'b11010011110010;
      12'b100010110001:
        _o_sv = 14'b11010011110111;
      12'b100010110010:
        _o_sv = 14'b11010011111101;
      12'b100010110011:
        _o_sv = 14'b11010100000011;
      12'b100010110100:
        _o_sv = 14'b11010100001000;
      12'b100010110101:
        _o_sv = 14'b11010100001110;
      12'b100010110110:
        _o_sv = 14'b11010100010100;
      12'b100010110111:
        _o_sv = 14'b11010100011010;
      12'b100010111000:
        _o_sv = 14'b11010100011111;
      12'b100010111001:
        _o_sv = 14'b11010100100101;
      12'b100010111010:
        _o_sv = 14'b11010100101011;
      12'b100010111011:
        _o_sv = 14'b11010100110000;
      12'b100010111100:
        _o_sv = 14'b11010100110110;
      12'b100010111101:
        _o_sv = 14'b11010100111100;
      12'b100010111110:
        _o_sv = 14'b11010101000010;
      12'b100010111111:
        _o_sv = 14'b11010101000111;
      12'b100011000000:
        _o_sv = 14'b11010101001101;
      12'b100011000001:
        _o_sv = 14'b11010101010011;
      12'b100011000010:
        _o_sv = 14'b11010101011000;
      12'b100011000011:
        _o_sv = 14'b11010101011110;
      12'b100011000100:
        _o_sv = 14'b11010101100100;
      12'b100011000101:
        _o_sv = 14'b11010101101010;
      12'b100011000110:
        _o_sv = 14'b11010101101111;
      12'b100011000111:
        _o_sv = 14'b11010101110101;
      12'b100011001000:
        _o_sv = 14'b11010101111011;
      12'b100011001001:
        _o_sv = 14'b11010110000000;
      12'b100011001010:
        _o_sv = 14'b11010110000110;
      12'b100011001011:
        _o_sv = 14'b11010110001100;
      12'b100011001100:
        _o_sv = 14'b11010110010010;
      12'b100011001101:
        _o_sv = 14'b11010110010111;
      12'b100011001110:
        _o_sv = 14'b11010110011101;
      12'b100011001111:
        _o_sv = 14'b11010110100011;
      12'b100011010000:
        _o_sv = 14'b11010110101000;
      12'b100011010001:
        _o_sv = 14'b11010110101110;
      12'b100011010010:
        _o_sv = 14'b11010110110100;
      12'b100011010011:
        _o_sv = 14'b11010110111010;
      12'b100011010100:
        _o_sv = 14'b11010110111111;
      12'b100011010101:
        _o_sv = 14'b11010111000101;
      12'b100011010110:
        _o_sv = 14'b11010111001011;
      12'b100011010111:
        _o_sv = 14'b11010111010000;
      12'b100011011000:
        _o_sv = 14'b11010111010110;
      12'b100011011001:
        _o_sv = 14'b11010111011100;
      12'b100011011010:
        _o_sv = 14'b11010111100001;
      12'b100011011011:
        _o_sv = 14'b11010111100111;
      12'b100011011100:
        _o_sv = 14'b11010111101101;
      12'b100011011101:
        _o_sv = 14'b11010111110011;
      12'b100011011110:
        _o_sv = 14'b11010111111000;
      12'b100011011111:
        _o_sv = 14'b11010111111110;
      12'b100011100000:
        _o_sv = 14'b11011000000100;
      12'b100011100001:
        _o_sv = 14'b11011000001001;
      12'b100011100010:
        _o_sv = 14'b11011000001111;
      12'b100011100011:
        _o_sv = 14'b11011000010101;
      12'b100011100100:
        _o_sv = 14'b11011000011010;
      12'b100011100101:
        _o_sv = 14'b11011000100000;
      12'b100011100110:
        _o_sv = 14'b11011000100110;
      12'b100011100111:
        _o_sv = 14'b11011000101011;
      12'b100011101000:
        _o_sv = 14'b11011000110001;
      12'b100011101001:
        _o_sv = 14'b11011000110111;
      12'b100011101010:
        _o_sv = 14'b11011000111101;
      12'b100011101011:
        _o_sv = 14'b11011001000010;
      12'b100011101100:
        _o_sv = 14'b11011001001000;
      12'b100011101101:
        _o_sv = 14'b11011001001110;
      12'b100011101110:
        _o_sv = 14'b11011001010011;
      12'b100011101111:
        _o_sv = 14'b11011001011001;
      12'b100011110000:
        _o_sv = 14'b11011001011111;
      12'b100011110001:
        _o_sv = 14'b11011001100100;
      12'b100011110010:
        _o_sv = 14'b11011001101010;
      12'b100011110011:
        _o_sv = 14'b11011001110000;
      12'b100011110100:
        _o_sv = 14'b11011001110101;
      12'b100011110101:
        _o_sv = 14'b11011001111011;
      12'b100011110110:
        _o_sv = 14'b11011010000001;
      12'b100011110111:
        _o_sv = 14'b11011010000110;
      12'b100011111000:
        _o_sv = 14'b11011010001100;
      12'b100011111001:
        _o_sv = 14'b11011010010010;
      12'b100011111010:
        _o_sv = 14'b11011010011000;
      12'b100011111011:
        _o_sv = 14'b11011010011101;
      12'b100011111100:
        _o_sv = 14'b11011010100011;
      12'b100011111101:
        _o_sv = 14'b11011010101001;
      12'b100011111110:
        _o_sv = 14'b11011010101110;
      12'b100011111111:
        _o_sv = 14'b11011010110100;
      12'b100100000000:
        _o_sv = 14'b11011010111010;
      12'b100100000001:
        _o_sv = 14'b11011010111111;
      12'b100100000010:
        _o_sv = 14'b11011011000101;
      12'b100100000011:
        _o_sv = 14'b11011011001011;
      12'b100100000100:
        _o_sv = 14'b11011011010000;
      12'b100100000101:
        _o_sv = 14'b11011011010110;
      12'b100100000110:
        _o_sv = 14'b11011011011100;
      12'b100100000111:
        _o_sv = 14'b11011011100001;
      12'b100100001000:
        _o_sv = 14'b11011011100111;
      12'b100100001001:
        _o_sv = 14'b11011011101101;
      12'b100100001010:
        _o_sv = 14'b11011011110010;
      12'b100100001011:
        _o_sv = 14'b11011011111000;
      12'b100100001100:
        _o_sv = 14'b11011011111110;
      12'b100100001101:
        _o_sv = 14'b11011100000011;
      12'b100100001110:
        _o_sv = 14'b11011100001001;
      12'b100100001111:
        _o_sv = 14'b11011100001111;
      12'b100100010000:
        _o_sv = 14'b11011100010100;
      12'b100100010001:
        _o_sv = 14'b11011100011010;
      12'b100100010010:
        _o_sv = 14'b11011100100000;
      12'b100100010011:
        _o_sv = 14'b11011100100101;
      12'b100100010100:
        _o_sv = 14'b11011100101011;
      12'b100100010101:
        _o_sv = 14'b11011100110001;
      12'b100100010110:
        _o_sv = 14'b11011100110110;
      12'b100100010111:
        _o_sv = 14'b11011100111100;
      12'b100100011000:
        _o_sv = 14'b11011101000010;
      12'b100100011001:
        _o_sv = 14'b11011101000111;
      12'b100100011010:
        _o_sv = 14'b11011101001101;
      12'b100100011011:
        _o_sv = 14'b11011101010011;
      12'b100100011100:
        _o_sv = 14'b11011101011000;
      12'b100100011101:
        _o_sv = 14'b11011101011110;
      12'b100100011110:
        _o_sv = 14'b11011101100100;
      12'b100100011111:
        _o_sv = 14'b11011101101001;
      12'b100100100000:
        _o_sv = 14'b11011101101111;
      12'b100100100001:
        _o_sv = 14'b11011101110101;
      12'b100100100010:
        _o_sv = 14'b11011101111010;
      12'b100100100011:
        _o_sv = 14'b11011110000000;
      12'b100100100100:
        _o_sv = 14'b11011110000110;
      12'b100100100101:
        _o_sv = 14'b11011110001011;
      12'b100100100110:
        _o_sv = 14'b11011110010001;
      12'b100100100111:
        _o_sv = 14'b11011110010111;
      12'b100100101000:
        _o_sv = 14'b11011110011100;
      12'b100100101001:
        _o_sv = 14'b11011110100010;
      12'b100100101010:
        _o_sv = 14'b11011110101000;
      12'b100100101011:
        _o_sv = 14'b11011110101101;
      12'b100100101100:
        _o_sv = 14'b11011110110011;
      12'b100100101101:
        _o_sv = 14'b11011110111001;
      12'b100100101110:
        _o_sv = 14'b11011110111110;
      12'b100100101111:
        _o_sv = 14'b11011111000100;
      12'b100100110000:
        _o_sv = 14'b11011111001010;
      12'b100100110001:
        _o_sv = 14'b11011111001111;
      12'b100100110010:
        _o_sv = 14'b11011111010101;
      12'b100100110011:
        _o_sv = 14'b11011111011011;
      12'b100100110100:
        _o_sv = 14'b11011111100000;
      12'b100100110101:
        _o_sv = 14'b11011111100110;
      12'b100100110110:
        _o_sv = 14'b11011111101100;
      12'b100100110111:
        _o_sv = 14'b11011111110001;
      12'b100100111000:
        _o_sv = 14'b11011111110111;
      12'b100100111001:
        _o_sv = 14'b11011111111101;
      12'b100100111010:
        _o_sv = 14'b11100000000010;
      12'b100100111011:
        _o_sv = 14'b11100000001000;
      12'b100100111100:
        _o_sv = 14'b11100000001101;
      12'b100100111101:
        _o_sv = 14'b11100000010011;
      12'b100100111110:
        _o_sv = 14'b11100000011001;
      12'b100100111111:
        _o_sv = 14'b11100000011110;
      12'b100101000000:
        _o_sv = 14'b11100000100100;
      12'b100101000001:
        _o_sv = 14'b11100000101010;
      12'b100101000010:
        _o_sv = 14'b11100000101111;
      12'b100101000011:
        _o_sv = 14'b11100000110101;
      12'b100101000100:
        _o_sv = 14'b11100000111011;
      12'b100101000101:
        _o_sv = 14'b11100001000000;
      12'b100101000110:
        _o_sv = 14'b11100001000110;
      12'b100101000111:
        _o_sv = 14'b11100001001100;
      12'b100101001000:
        _o_sv = 14'b11100001010001;
      12'b100101001001:
        _o_sv = 14'b11100001010111;
      12'b100101001010:
        _o_sv = 14'b11100001011101;
      12'b100101001011:
        _o_sv = 14'b11100001100010;
      12'b100101001100:
        _o_sv = 14'b11100001101000;
      12'b100101001101:
        _o_sv = 14'b11100001101101;
      12'b100101001110:
        _o_sv = 14'b11100001110011;
      12'b100101001111:
        _o_sv = 14'b11100001111001;
      12'b100101010000:
        _o_sv = 14'b11100001111110;
      12'b100101010001:
        _o_sv = 14'b11100010000100;
      12'b100101010010:
        _o_sv = 14'b11100010001010;
      12'b100101010011:
        _o_sv = 14'b11100010001111;
      12'b100101010100:
        _o_sv = 14'b11100010010101;
      12'b100101010101:
        _o_sv = 14'b11100010011011;
      12'b100101010110:
        _o_sv = 14'b11100010100000;
      12'b100101010111:
        _o_sv = 14'b11100010100110;
      12'b100101011000:
        _o_sv = 14'b11100010101011;
      12'b100101011001:
        _o_sv = 14'b11100010110001;
      12'b100101011010:
        _o_sv = 14'b11100010110111;
      12'b100101011011:
        _o_sv = 14'b11100010111100;
      12'b100101011100:
        _o_sv = 14'b11100011000010;
      12'b100101011101:
        _o_sv = 14'b11100011001000;
      12'b100101011110:
        _o_sv = 14'b11100011001101;
      12'b100101011111:
        _o_sv = 14'b11100011010011;
      12'b100101100000:
        _o_sv = 14'b11100011011000;
      12'b100101100001:
        _o_sv = 14'b11100011011110;
      12'b100101100010:
        _o_sv = 14'b11100011100100;
      12'b100101100011:
        _o_sv = 14'b11100011101001;
      12'b100101100100:
        _o_sv = 14'b11100011101111;
      12'b100101100101:
        _o_sv = 14'b11100011110101;
      12'b100101100110:
        _o_sv = 14'b11100011111010;
      12'b100101100111:
        _o_sv = 14'b11100100000000;
      12'b100101101000:
        _o_sv = 14'b11100100000110;
      12'b100101101001:
        _o_sv = 14'b11100100001011;
      12'b100101101010:
        _o_sv = 14'b11100100010001;
      12'b100101101011:
        _o_sv = 14'b11100100010110;
      12'b100101101100:
        _o_sv = 14'b11100100011100;
      12'b100101101101:
        _o_sv = 14'b11100100100010;
      12'b100101101110:
        _o_sv = 14'b11100100100111;
      12'b100101101111:
        _o_sv = 14'b11100100101101;
      12'b100101110000:
        _o_sv = 14'b11100100110010;
      12'b100101110001:
        _o_sv = 14'b11100100111000;
      12'b100101110010:
        _o_sv = 14'b11100100111110;
      12'b100101110011:
        _o_sv = 14'b11100101000011;
      12'b100101110100:
        _o_sv = 14'b11100101001001;
      12'b100101110101:
        _o_sv = 14'b11100101001111;
      12'b100101110110:
        _o_sv = 14'b11100101010100;
      12'b100101110111:
        _o_sv = 14'b11100101011010;
      12'b100101111000:
        _o_sv = 14'b11100101011111;
      12'b100101111001:
        _o_sv = 14'b11100101100101;
      12'b100101111010:
        _o_sv = 14'b11100101101011;
      12'b100101111011:
        _o_sv = 14'b11100101110000;
      12'b100101111100:
        _o_sv = 14'b11100101110110;
      12'b100101111101:
        _o_sv = 14'b11100101111100;
      12'b100101111110:
        _o_sv = 14'b11100110000001;
      12'b100101111111:
        _o_sv = 14'b11100110000111;
      12'b100110000000:
        _o_sv = 14'b11100110001100;
      12'b100110000001:
        _o_sv = 14'b11100110010010;
      12'b100110000010:
        _o_sv = 14'b11100110011000;
      12'b100110000011:
        _o_sv = 14'b11100110011101;
      12'b100110000100:
        _o_sv = 14'b11100110100011;
      12'b100110000101:
        _o_sv = 14'b11100110101000;
      12'b100110000110:
        _o_sv = 14'b11100110101110;
      12'b100110000111:
        _o_sv = 14'b11100110110100;
      12'b100110001000:
        _o_sv = 14'b11100110111001;
      12'b100110001001:
        _o_sv = 14'b11100110111111;
      12'b100110001010:
        _o_sv = 14'b11100111000100;
      12'b100110001011:
        _o_sv = 14'b11100111001010;
      12'b100110001100:
        _o_sv = 14'b11100111010000;
      12'b100110001101:
        _o_sv = 14'b11100111010101;
      12'b100110001110:
        _o_sv = 14'b11100111011011;
      12'b100110001111:
        _o_sv = 14'b11100111100000;
      12'b100110010000:
        _o_sv = 14'b11100111100110;
      12'b100110010001:
        _o_sv = 14'b11100111101100;
      12'b100110010010:
        _o_sv = 14'b11100111110001;
      12'b100110010011:
        _o_sv = 14'b11100111110111;
      12'b100110010100:
        _o_sv = 14'b11100111111101;
      12'b100110010101:
        _o_sv = 14'b11101000000010;
      12'b100110010110:
        _o_sv = 14'b11101000001000;
      12'b100110010111:
        _o_sv = 14'b11101000001101;
      12'b100110011000:
        _o_sv = 14'b11101000010011;
      12'b100110011001:
        _o_sv = 14'b11101000011001;
      12'b100110011010:
        _o_sv = 14'b11101000011110;
      12'b100110011011:
        _o_sv = 14'b11101000100100;
      12'b100110011100:
        _o_sv = 14'b11101000101001;
      12'b100110011101:
        _o_sv = 14'b11101000101111;
      12'b100110011110:
        _o_sv = 14'b11101000110100;
      12'b100110011111:
        _o_sv = 14'b11101000111010;
      12'b100110100000:
        _o_sv = 14'b11101001000000;
      12'b100110100001:
        _o_sv = 14'b11101001000101;
      12'b100110100010:
        _o_sv = 14'b11101001001011;
      12'b100110100011:
        _o_sv = 14'b11101001010000;
      12'b100110100100:
        _o_sv = 14'b11101001010110;
      12'b100110100101:
        _o_sv = 14'b11101001011100;
      12'b100110100110:
        _o_sv = 14'b11101001100001;
      12'b100110100111:
        _o_sv = 14'b11101001100111;
      12'b100110101000:
        _o_sv = 14'b11101001101100;
      12'b100110101001:
        _o_sv = 14'b11101001110010;
      12'b100110101010:
        _o_sv = 14'b11101001111000;
      12'b100110101011:
        _o_sv = 14'b11101001111101;
      12'b100110101100:
        _o_sv = 14'b11101010000011;
      12'b100110101101:
        _o_sv = 14'b11101010001000;
      12'b100110101110:
        _o_sv = 14'b11101010001110;
      12'b100110101111:
        _o_sv = 14'b11101010010100;
      12'b100110110000:
        _o_sv = 14'b11101010011001;
      12'b100110110001:
        _o_sv = 14'b11101010011111;
      12'b100110110010:
        _o_sv = 14'b11101010100100;
      12'b100110110011:
        _o_sv = 14'b11101010101010;
      12'b100110110100:
        _o_sv = 14'b11101010101111;
      12'b100110110101:
        _o_sv = 14'b11101010110101;
      12'b100110110110:
        _o_sv = 14'b11101010111011;
      12'b100110110111:
        _o_sv = 14'b11101011000000;
      12'b100110111000:
        _o_sv = 14'b11101011000110;
      12'b100110111001:
        _o_sv = 14'b11101011001011;
      12'b100110111010:
        _o_sv = 14'b11101011010001;
      12'b100110111011:
        _o_sv = 14'b11101011010111;
      12'b100110111100:
        _o_sv = 14'b11101011011100;
      12'b100110111101:
        _o_sv = 14'b11101011100010;
      12'b100110111110:
        _o_sv = 14'b11101011100111;
      12'b100110111111:
        _o_sv = 14'b11101011101101;
      12'b100111000000:
        _o_sv = 14'b11101011110010;
      12'b100111000001:
        _o_sv = 14'b11101011111000;
      12'b100111000010:
        _o_sv = 14'b11101011111110;
      12'b100111000011:
        _o_sv = 14'b11101100000011;
      12'b100111000100:
        _o_sv = 14'b11101100001001;
      12'b100111000101:
        _o_sv = 14'b11101100001110;
      12'b100111000110:
        _o_sv = 14'b11101100010100;
      12'b100111000111:
        _o_sv = 14'b11101100011001;
      12'b100111001000:
        _o_sv = 14'b11101100011111;
      12'b100111001001:
        _o_sv = 14'b11101100100101;
      12'b100111001010:
        _o_sv = 14'b11101100101010;
      12'b100111001011:
        _o_sv = 14'b11101100110000;
      12'b100111001100:
        _o_sv = 14'b11101100110101;
      12'b100111001101:
        _o_sv = 14'b11101100111011;
      12'b100111001110:
        _o_sv = 14'b11101101000000;
      12'b100111001111:
        _o_sv = 14'b11101101000110;
      12'b100111010000:
        _o_sv = 14'b11101101001100;
      12'b100111010001:
        _o_sv = 14'b11101101010001;
      12'b100111010010:
        _o_sv = 14'b11101101010111;
      12'b100111010011:
        _o_sv = 14'b11101101011100;
      12'b100111010100:
        _o_sv = 14'b11101101100010;
      12'b100111010101:
        _o_sv = 14'b11101101100111;
      12'b100111010110:
        _o_sv = 14'b11101101101101;
      12'b100111010111:
        _o_sv = 14'b11101101110011;
      12'b100111011000:
        _o_sv = 14'b11101101111000;
      12'b100111011001:
        _o_sv = 14'b11101101111110;
      12'b100111011010:
        _o_sv = 14'b11101110000011;
      12'b100111011011:
        _o_sv = 14'b11101110001001;
      12'b100111011100:
        _o_sv = 14'b11101110001110;
      12'b100111011101:
        _o_sv = 14'b11101110010100;
      12'b100111011110:
        _o_sv = 14'b11101110011001;
      12'b100111011111:
        _o_sv = 14'b11101110011111;
      12'b100111100000:
        _o_sv = 14'b11101110100101;
      12'b100111100001:
        _o_sv = 14'b11101110101010;
      12'b100111100010:
        _o_sv = 14'b11101110110000;
      12'b100111100011:
        _o_sv = 14'b11101110110101;
      12'b100111100100:
        _o_sv = 14'b11101110111011;
      12'b100111100101:
        _o_sv = 14'b11101111000000;
      12'b100111100110:
        _o_sv = 14'b11101111000110;
      12'b100111100111:
        _o_sv = 14'b11101111001100;
      12'b100111101000:
        _o_sv = 14'b11101111010001;
      12'b100111101001:
        _o_sv = 14'b11101111010111;
      12'b100111101010:
        _o_sv = 14'b11101111011100;
      12'b100111101011:
        _o_sv = 14'b11101111100010;
      12'b100111101100:
        _o_sv = 14'b11101111100111;
      12'b100111101101:
        _o_sv = 14'b11101111101101;
      12'b100111101110:
        _o_sv = 14'b11101111110010;
      12'b100111101111:
        _o_sv = 14'b11101111111000;
      12'b100111110000:
        _o_sv = 14'b11101111111101;
      12'b100111110001:
        _o_sv = 14'b11110000000011;
      12'b100111110010:
        _o_sv = 14'b11110000001001;
      12'b100111110011:
        _o_sv = 14'b11110000001110;
      12'b100111110100:
        _o_sv = 14'b11110000010100;
      12'b100111110101:
        _o_sv = 14'b11110000011001;
      12'b100111110110:
        _o_sv = 14'b11110000011111;
      12'b100111110111:
        _o_sv = 14'b11110000100100;
      12'b100111111000:
        _o_sv = 14'b11110000101010;
      12'b100111111001:
        _o_sv = 14'b11110000101111;
      12'b100111111010:
        _o_sv = 14'b11110000110101;
      12'b100111111011:
        _o_sv = 14'b11110000111011;
      12'b100111111100:
        _o_sv = 14'b11110001000000;
      12'b100111111101:
        _o_sv = 14'b11110001000110;
      12'b100111111110:
        _o_sv = 14'b11110001001011;
      12'b100111111111:
        _o_sv = 14'b11110001010001;
      12'b101000000000:
        _o_sv = 14'b11110001010110;
      12'b101000000001:
        _o_sv = 14'b11110001011100;
      12'b101000000010:
        _o_sv = 14'b11110001100001;
      12'b101000000011:
        _o_sv = 14'b11110001100111;
      12'b101000000100:
        _o_sv = 14'b11110001101100;
      12'b101000000101:
        _o_sv = 14'b11110001110010;
      12'b101000000110:
        _o_sv = 14'b11110001110111;
      12'b101000000111:
        _o_sv = 14'b11110001111101;
      12'b101000001000:
        _o_sv = 14'b11110010000011;
      12'b101000001001:
        _o_sv = 14'b11110010001000;
      12'b101000001010:
        _o_sv = 14'b11110010001110;
      12'b101000001011:
        _o_sv = 14'b11110010010011;
      12'b101000001100:
        _o_sv = 14'b11110010011001;
      12'b101000001101:
        _o_sv = 14'b11110010011110;
      12'b101000001110:
        _o_sv = 14'b11110010100100;
      12'b101000001111:
        _o_sv = 14'b11110010101001;
      12'b101000010000:
        _o_sv = 14'b11110010101111;
      12'b101000010001:
        _o_sv = 14'b11110010110100;
      12'b101000010010:
        _o_sv = 14'b11110010111010;
      12'b101000010011:
        _o_sv = 14'b11110010111111;
      12'b101000010100:
        _o_sv = 14'b11110011000101;
      12'b101000010101:
        _o_sv = 14'b11110011001010;
      12'b101000010110:
        _o_sv = 14'b11110011010000;
      12'b101000010111:
        _o_sv = 14'b11110011010110;
      12'b101000011000:
        _o_sv = 14'b11110011011011;
      12'b101000011001:
        _o_sv = 14'b11110011100001;
      12'b101000011010:
        _o_sv = 14'b11110011100110;
      12'b101000011011:
        _o_sv = 14'b11110011101100;
      12'b101000011100:
        _o_sv = 14'b11110011110001;
      12'b101000011101:
        _o_sv = 14'b11110011110111;
      12'b101000011110:
        _o_sv = 14'b11110011111100;
      12'b101000011111:
        _o_sv = 14'b11110100000010;
      12'b101000100000:
        _o_sv = 14'b11110100000111;
      12'b101000100001:
        _o_sv = 14'b11110100001101;
      12'b101000100010:
        _o_sv = 14'b11110100010010;
      12'b101000100011:
        _o_sv = 14'b11110100011000;
      12'b101000100100:
        _o_sv = 14'b11110100011101;
      12'b101000100101:
        _o_sv = 14'b11110100100011;
      12'b101000100110:
        _o_sv = 14'b11110100101000;
      12'b101000100111:
        _o_sv = 14'b11110100101110;
      12'b101000101000:
        _o_sv = 14'b11110100110011;
      12'b101000101001:
        _o_sv = 14'b11110100111001;
      12'b101000101010:
        _o_sv = 14'b11110100111110;
      12'b101000101011:
        _o_sv = 14'b11110101000100;
      12'b101000101100:
        _o_sv = 14'b11110101001001;
      12'b101000101101:
        _o_sv = 14'b11110101001111;
      12'b101000101110:
        _o_sv = 14'b11110101010101;
      12'b101000101111:
        _o_sv = 14'b11110101011010;
      12'b101000110000:
        _o_sv = 14'b11110101100000;
      12'b101000110001:
        _o_sv = 14'b11110101100101;
      12'b101000110010:
        _o_sv = 14'b11110101101011;
      12'b101000110011:
        _o_sv = 14'b11110101110000;
      12'b101000110100:
        _o_sv = 14'b11110101110110;
      12'b101000110101:
        _o_sv = 14'b11110101111011;
      12'b101000110110:
        _o_sv = 14'b11110110000001;
      12'b101000110111:
        _o_sv = 14'b11110110000110;
      12'b101000111000:
        _o_sv = 14'b11110110001100;
      12'b101000111001:
        _o_sv = 14'b11110110010001;
      12'b101000111010:
        _o_sv = 14'b11110110010111;
      12'b101000111011:
        _o_sv = 14'b11110110011100;
      12'b101000111100:
        _o_sv = 14'b11110110100010;
      12'b101000111101:
        _o_sv = 14'b11110110100111;
      12'b101000111110:
        _o_sv = 14'b11110110101101;
      12'b101000111111:
        _o_sv = 14'b11110110110010;
      12'b101001000000:
        _o_sv = 14'b11110110111000;
      12'b101001000001:
        _o_sv = 14'b11110110111101;
      12'b101001000010:
        _o_sv = 14'b11110111000011;
      12'b101001000011:
        _o_sv = 14'b11110111001000;
      12'b101001000100:
        _o_sv = 14'b11110111001110;
      12'b101001000101:
        _o_sv = 14'b11110111010011;
      12'b101001000110:
        _o_sv = 14'b11110111011001;
      12'b101001000111:
        _o_sv = 14'b11110111011110;
      12'b101001001000:
        _o_sv = 14'b11110111100100;
      12'b101001001001:
        _o_sv = 14'b11110111101001;
      12'b101001001010:
        _o_sv = 14'b11110111101111;
      12'b101001001011:
        _o_sv = 14'b11110111110100;
      12'b101001001100:
        _o_sv = 14'b11110111111010;
      12'b101001001101:
        _o_sv = 14'b11110111111111;
      12'b101001001110:
        _o_sv = 14'b11111000000101;
      12'b101001001111:
        _o_sv = 14'b11111000001010;
      12'b101001010000:
        _o_sv = 14'b11111000010000;
      12'b101001010001:
        _o_sv = 14'b11111000010101;
      12'b101001010010:
        _o_sv = 14'b11111000011011;
      12'b101001010011:
        _o_sv = 14'b11111000100000;
      12'b101001010100:
        _o_sv = 14'b11111000100110;
      12'b101001010101:
        _o_sv = 14'b11111000101011;
      12'b101001010110:
        _o_sv = 14'b11111000110001;
      12'b101001010111:
        _o_sv = 14'b11111000110110;
      12'b101001011000:
        _o_sv = 14'b11111000111100;
      12'b101001011001:
        _o_sv = 14'b11111001000001;
      12'b101001011010:
        _o_sv = 14'b11111001000111;
      12'b101001011011:
        _o_sv = 14'b11111001001100;
      12'b101001011100:
        _o_sv = 14'b11111001010010;
      12'b101001011101:
        _o_sv = 14'b11111001010111;
      12'b101001011110:
        _o_sv = 14'b11111001011101;
      12'b101001011111:
        _o_sv = 14'b11111001100010;
      12'b101001100000:
        _o_sv = 14'b11111001101000;
      12'b101001100001:
        _o_sv = 14'b11111001101101;
      12'b101001100010:
        _o_sv = 14'b11111001110011;
      12'b101001100011:
        _o_sv = 14'b11111001111000;
      12'b101001100100:
        _o_sv = 14'b11111001111101;
      12'b101001100101:
        _o_sv = 14'b11111010000011;
      12'b101001100110:
        _o_sv = 14'b11111010001000;
      12'b101001100111:
        _o_sv = 14'b11111010001110;
      12'b101001101000:
        _o_sv = 14'b11111010010011;
      12'b101001101001:
        _o_sv = 14'b11111010011001;
      12'b101001101010:
        _o_sv = 14'b11111010011110;
      12'b101001101011:
        _o_sv = 14'b11111010100100;
      12'b101001101100:
        _o_sv = 14'b11111010101001;
      12'b101001101101:
        _o_sv = 14'b11111010101111;
      12'b101001101110:
        _o_sv = 14'b11111010110100;
      12'b101001101111:
        _o_sv = 14'b11111010111010;
      12'b101001110000:
        _o_sv = 14'b11111010111111;
      12'b101001110001:
        _o_sv = 14'b11111011000101;
      12'b101001110010:
        _o_sv = 14'b11111011001010;
      12'b101001110011:
        _o_sv = 14'b11111011010000;
      12'b101001110100:
        _o_sv = 14'b11111011010101;
      12'b101001110101:
        _o_sv = 14'b11111011011011;
      12'b101001110110:
        _o_sv = 14'b11111011100000;
      12'b101001110111:
        _o_sv = 14'b11111011100110;
      12'b101001111000:
        _o_sv = 14'b11111011101011;
      12'b101001111001:
        _o_sv = 14'b11111011110001;
      12'b101001111010:
        _o_sv = 14'b11111011110110;
      12'b101001111011:
        _o_sv = 14'b11111011111011;
      12'b101001111100:
        _o_sv = 14'b11111100000001;
      12'b101001111101:
        _o_sv = 14'b11111100000110;
      12'b101001111110:
        _o_sv = 14'b11111100001100;
      12'b101001111111:
        _o_sv = 14'b11111100010001;
      12'b101010000000:
        _o_sv = 14'b11111100010111;
      12'b101010000001:
        _o_sv = 14'b11111100011100;
      12'b101010000010:
        _o_sv = 14'b11111100100010;
      12'b101010000011:
        _o_sv = 14'b11111100100111;
      12'b101010000100:
        _o_sv = 14'b11111100101101;
      12'b101010000101:
        _o_sv = 14'b11111100110010;
      12'b101010000110:
        _o_sv = 14'b11111100111000;
      12'b101010000111:
        _o_sv = 14'b11111100111101;
      12'b101010001000:
        _o_sv = 14'b11111101000011;
      12'b101010001001:
        _o_sv = 14'b11111101001000;
      12'b101010001010:
        _o_sv = 14'b11111101001101;
      12'b101010001011:
        _o_sv = 14'b11111101010011;
      12'b101010001100:
        _o_sv = 14'b11111101011000;
      12'b101010001101:
        _o_sv = 14'b11111101011110;
      12'b101010001110:
        _o_sv = 14'b11111101100011;
      12'b101010001111:
        _o_sv = 14'b11111101101001;
      12'b101010010000:
        _o_sv = 14'b11111101101110;
      12'b101010010001:
        _o_sv = 14'b11111101110100;
      12'b101010010010:
        _o_sv = 14'b11111101111001;
      12'b101010010011:
        _o_sv = 14'b11111101111111;
      12'b101010010100:
        _o_sv = 14'b11111110000100;
      12'b101010010101:
        _o_sv = 14'b11111110001001;
      12'b101010010110:
        _o_sv = 14'b11111110001111;
      12'b101010010111:
        _o_sv = 14'b11111110010100;
      12'b101010011000:
        _o_sv = 14'b11111110011010;
      12'b101010011001:
        _o_sv = 14'b11111110011111;
      12'b101010011010:
        _o_sv = 14'b11111110100101;
      12'b101010011011:
        _o_sv = 14'b11111110101010;
      12'b101010011100:
        _o_sv = 14'b11111110110000;
      12'b101010011101:
        _o_sv = 14'b11111110110101;
      12'b101010011110:
        _o_sv = 14'b11111110111011;
      12'b101010011111:
        _o_sv = 14'b11111111000000;
      12'b101010100000:
        _o_sv = 14'b11111111000101;
      12'b101010100001:
        _o_sv = 14'b11111111001011;
      12'b101010100010:
        _o_sv = 14'b11111111010000;
      12'b101010100011:
        _o_sv = 14'b11111111010110;
      12'b101010100100:
        _o_sv = 14'b11111111011011;
      12'b101010100101:
        _o_sv = 14'b11111111100001;
      12'b101010100110:
        _o_sv = 14'b11111111100110;
      12'b101010100111:
        _o_sv = 14'b11111111101100;
      12'b101010101000:
        _o_sv = 14'b11111111110001;
      12'b101010101001:
        _o_sv = 14'b11111111110110;
      12'b101010101010:
        _o_sv = 14'b11111111111100;
      12'b101010101011:
        _o_sv = 15'b100000000000001;
      12'b101010101100:
        _o_sv = 15'b100000000000111;
      12'b101010101101:
        _o_sv = 15'b100000000001100;
      12'b101010101110:
        _o_sv = 15'b100000000010010;
      12'b101010101111:
        _o_sv = 15'b100000000010111;
      12'b101010110000:
        _o_sv = 15'b100000000011101;
      12'b101010110001:
        _o_sv = 15'b100000000100010;
      12'b101010110010:
        _o_sv = 15'b100000000100111;
      12'b101010110011:
        _o_sv = 15'b100000000101101;
      12'b101010110100:
        _o_sv = 15'b100000000110010;
      12'b101010110101:
        _o_sv = 15'b100000000111000;
      12'b101010110110:
        _o_sv = 15'b100000000111101;
      12'b101010110111:
        _o_sv = 15'b100000001000011;
      12'b101010111000:
        _o_sv = 15'b100000001001000;
      12'b101010111001:
        _o_sv = 15'b100000001001101;
      12'b101010111010:
        _o_sv = 15'b100000001010011;
      12'b101010111011:
        _o_sv = 15'b100000001011000;
      12'b101010111100:
        _o_sv = 15'b100000001011110;
      12'b101010111101:
        _o_sv = 15'b100000001100011;
      12'b101010111110:
        _o_sv = 15'b100000001101001;
      12'b101010111111:
        _o_sv = 15'b100000001101110;
      12'b101011000000:
        _o_sv = 15'b100000001110011;
      12'b101011000001:
        _o_sv = 15'b100000001111001;
      12'b101011000010:
        _o_sv = 15'b100000001111110;
      12'b101011000011:
        _o_sv = 15'b100000010000100;
      12'b101011000100:
        _o_sv = 15'b100000010001001;
      12'b101011000101:
        _o_sv = 15'b100000010001111;
      12'b101011000110:
        _o_sv = 15'b100000010010100;
      12'b101011000111:
        _o_sv = 15'b100000010011001;
      12'b101011001000:
        _o_sv = 15'b100000010011111;
      12'b101011001001:
        _o_sv = 15'b100000010100100;
      12'b101011001010:
        _o_sv = 15'b100000010101010;
      12'b101011001011:
        _o_sv = 15'b100000010101111;
      12'b101011001100:
        _o_sv = 15'b100000010110101;
      12'b101011001101:
        _o_sv = 15'b100000010111010;
      12'b101011001110:
        _o_sv = 15'b100000010111111;
      12'b101011001111:
        _o_sv = 15'b100000011000101;
      12'b101011010000:
        _o_sv = 15'b100000011001010;
      12'b101011010001:
        _o_sv = 15'b100000011010000;
      12'b101011010010:
        _o_sv = 15'b100000011010101;
      12'b101011010011:
        _o_sv = 15'b100000011011010;
      12'b101011010100:
        _o_sv = 15'b100000011100000;
      12'b101011010101:
        _o_sv = 15'b100000011100101;
      12'b101011010110:
        _o_sv = 15'b100000011101011;
      12'b101011010111:
        _o_sv = 15'b100000011110000;
      12'b101011011000:
        _o_sv = 15'b100000011110110;
      12'b101011011001:
        _o_sv = 15'b100000011111011;
      12'b101011011010:
        _o_sv = 15'b100000100000000;
      12'b101011011011:
        _o_sv = 15'b100000100000110;
      12'b101011011100:
        _o_sv = 15'b100000100001011;
      12'b101011011101:
        _o_sv = 15'b100000100010001;
      12'b101011011110:
        _o_sv = 15'b100000100010110;
      12'b101011011111:
        _o_sv = 15'b100000100011011;
      12'b101011100000:
        _o_sv = 15'b100000100100001;
      12'b101011100001:
        _o_sv = 15'b100000100100110;
      12'b101011100010:
        _o_sv = 15'b100000100101100;
      12'b101011100011:
        _o_sv = 15'b100000100110001;
      12'b101011100100:
        _o_sv = 15'b100000100110110;
      12'b101011100101:
        _o_sv = 15'b100000100111100;
      12'b101011100110:
        _o_sv = 15'b100000101000001;
      12'b101011100111:
        _o_sv = 15'b100000101000111;
      12'b101011101000:
        _o_sv = 15'b100000101001100;
      12'b101011101001:
        _o_sv = 15'b100000101010010;
      12'b101011101010:
        _o_sv = 15'b100000101010111;
      12'b101011101011:
        _o_sv = 15'b100000101011100;
      12'b101011101100:
        _o_sv = 15'b100000101100010;
      12'b101011101101:
        _o_sv = 15'b100000101100111;
      12'b101011101110:
        _o_sv = 15'b100000101101101;
      12'b101011101111:
        _o_sv = 15'b100000101110010;
      12'b101011110000:
        _o_sv = 15'b100000101110111;
      12'b101011110001:
        _o_sv = 15'b100000101111101;
      12'b101011110010:
        _o_sv = 15'b100000110000010;
      12'b101011110011:
        _o_sv = 15'b100000110001000;
      12'b101011110100:
        _o_sv = 15'b100000110001101;
      12'b101011110101:
        _o_sv = 15'b100000110010010;
      12'b101011110110:
        _o_sv = 15'b100000110011000;
      12'b101011110111:
        _o_sv = 15'b100000110011101;
      12'b101011111000:
        _o_sv = 15'b100000110100010;
      12'b101011111001:
        _o_sv = 15'b100000110101000;
      12'b101011111010:
        _o_sv = 15'b100000110101101;
      12'b101011111011:
        _o_sv = 15'b100000110110011;
      12'b101011111100:
        _o_sv = 15'b100000110111000;
      12'b101011111101:
        _o_sv = 15'b100000110111101;
      12'b101011111110:
        _o_sv = 15'b100000111000011;
      12'b101011111111:
        _o_sv = 15'b100000111001000;
      12'b101100000000:
        _o_sv = 15'b100000111001110;
      12'b101100000001:
        _o_sv = 15'b100000111010011;
      12'b101100000010:
        _o_sv = 15'b100000111011000;
      12'b101100000011:
        _o_sv = 15'b100000111011110;
      12'b101100000100:
        _o_sv = 15'b100000111100011;
      12'b101100000101:
        _o_sv = 15'b100000111101001;
      12'b101100000110:
        _o_sv = 15'b100000111101110;
      12'b101100000111:
        _o_sv = 15'b100000111110011;
      12'b101100001000:
        _o_sv = 15'b100000111111001;
      12'b101100001001:
        _o_sv = 15'b100000111111110;
      12'b101100001010:
        _o_sv = 15'b100001000000011;
      12'b101100001011:
        _o_sv = 15'b100001000001001;
      12'b101100001100:
        _o_sv = 15'b100001000001110;
      12'b101100001101:
        _o_sv = 15'b100001000010100;
      12'b101100001110:
        _o_sv = 15'b100001000011001;
      12'b101100001111:
        _o_sv = 15'b100001000011110;
      12'b101100010000:
        _o_sv = 15'b100001000100100;
      12'b101100010001:
        _o_sv = 15'b100001000101001;
      12'b101100010010:
        _o_sv = 15'b100001000101111;
      12'b101100010011:
        _o_sv = 15'b100001000110100;
      12'b101100010100:
        _o_sv = 15'b100001000111001;
      12'b101100010101:
        _o_sv = 15'b100001000111111;
      12'b101100010110:
        _o_sv = 15'b100001001000100;
      12'b101100010111:
        _o_sv = 15'b100001001001001;
      12'b101100011000:
        _o_sv = 15'b100001001001111;
      12'b101100011001:
        _o_sv = 15'b100001001010100;
      12'b101100011010:
        _o_sv = 15'b100001001011010;
      12'b101100011011:
        _o_sv = 15'b100001001011111;
      12'b101100011100:
        _o_sv = 15'b100001001100100;
      12'b101100011101:
        _o_sv = 15'b100001001101010;
      12'b101100011110:
        _o_sv = 15'b100001001101111;
      12'b101100011111:
        _o_sv = 15'b100001001110100;
      12'b101100100000:
        _o_sv = 15'b100001001111010;
      12'b101100100001:
        _o_sv = 15'b100001001111111;
      12'b101100100010:
        _o_sv = 15'b100001010000100;
      12'b101100100011:
        _o_sv = 15'b100001010001010;
      12'b101100100100:
        _o_sv = 15'b100001010001111;
      12'b101100100101:
        _o_sv = 15'b100001010010101;
      12'b101100100110:
        _o_sv = 15'b100001010011010;
      12'b101100100111:
        _o_sv = 15'b100001010011111;
      12'b101100101000:
        _o_sv = 15'b100001010100101;
      12'b101100101001:
        _o_sv = 15'b100001010101010;
      12'b101100101010:
        _o_sv = 15'b100001010101111;
      12'b101100101011:
        _o_sv = 15'b100001010110101;
      12'b101100101100:
        _o_sv = 15'b100001010111010;
      12'b101100101101:
        _o_sv = 15'b100001011000000;
      12'b101100101110:
        _o_sv = 15'b100001011000101;
      12'b101100101111:
        _o_sv = 15'b100001011001010;
      12'b101100110000:
        _o_sv = 15'b100001011010000;
      12'b101100110001:
        _o_sv = 15'b100001011010101;
      12'b101100110010:
        _o_sv = 15'b100001011011010;
      12'b101100110011:
        _o_sv = 15'b100001011100000;
      12'b101100110100:
        _o_sv = 15'b100001011100101;
      12'b101100110101:
        _o_sv = 15'b100001011101010;
      12'b101100110110:
        _o_sv = 15'b100001011110000;
      12'b101100110111:
        _o_sv = 15'b100001011110101;
      12'b101100111000:
        _o_sv = 15'b100001011111010;
      12'b101100111001:
        _o_sv = 15'b100001100000000;
      12'b101100111010:
        _o_sv = 15'b100001100000101;
      12'b101100111011:
        _o_sv = 15'b100001100001011;
      12'b101100111100:
        _o_sv = 15'b100001100010000;
      12'b101100111101:
        _o_sv = 15'b100001100010101;
      12'b101100111110:
        _o_sv = 15'b100001100011011;
      12'b101100111111:
        _o_sv = 15'b100001100100000;
      12'b101101000000:
        _o_sv = 15'b100001100100101;
      12'b101101000001:
        _o_sv = 15'b100001100101011;
      12'b101101000010:
        _o_sv = 15'b100001100110000;
      12'b101101000011:
        _o_sv = 15'b100001100110101;
      12'b101101000100:
        _o_sv = 15'b100001100111011;
      12'b101101000101:
        _o_sv = 15'b100001101000000;
      12'b101101000110:
        _o_sv = 15'b100001101000101;
      12'b101101000111:
        _o_sv = 15'b100001101001011;
      12'b101101001000:
        _o_sv = 15'b100001101010000;
      12'b101101001001:
        _o_sv = 15'b100001101010101;
      12'b101101001010:
        _o_sv = 15'b100001101011011;
      12'b101101001011:
        _o_sv = 15'b100001101100000;
      12'b101101001100:
        _o_sv = 15'b100001101100101;
      12'b101101001101:
        _o_sv = 15'b100001101101011;
      12'b101101001110:
        _o_sv = 15'b100001101110000;
      12'b101101001111:
        _o_sv = 15'b100001101110101;
      12'b101101010000:
        _o_sv = 15'b100001101111011;
      12'b101101010001:
        _o_sv = 15'b100001110000000;
      12'b101101010010:
        _o_sv = 15'b100001110000101;
      12'b101101010011:
        _o_sv = 15'b100001110001011;
      12'b101101010100:
        _o_sv = 15'b100001110010000;
      12'b101101010101:
        _o_sv = 15'b100001110010101;
      12'b101101010110:
        _o_sv = 15'b100001110011011;
      12'b101101010111:
        _o_sv = 15'b100001110100000;
      12'b101101011000:
        _o_sv = 15'b100001110100101;
      12'b101101011001:
        _o_sv = 15'b100001110101011;
      12'b101101011010:
        _o_sv = 15'b100001110110000;
      12'b101101011011:
        _o_sv = 15'b100001110110101;
      12'b101101011100:
        _o_sv = 15'b100001110111011;
      12'b101101011101:
        _o_sv = 15'b100001111000000;
      12'b101101011110:
        _o_sv = 15'b100001111000101;
      12'b101101011111:
        _o_sv = 15'b100001111001011;
      12'b101101100000:
        _o_sv = 15'b100001111010000;
      12'b101101100001:
        _o_sv = 15'b100001111010101;
      12'b101101100010:
        _o_sv = 15'b100001111011011;
      12'b101101100011:
        _o_sv = 15'b100001111100000;
      12'b101101100100:
        _o_sv = 15'b100001111100101;
      12'b101101100101:
        _o_sv = 15'b100001111101011;
      12'b101101100110:
        _o_sv = 15'b100001111110000;
      12'b101101100111:
        _o_sv = 15'b100001111110101;
      12'b101101101000:
        _o_sv = 15'b100001111111011;
      12'b101101101001:
        _o_sv = 15'b100010000000000;
      12'b101101101010:
        _o_sv = 15'b100010000000101;
      12'b101101101011:
        _o_sv = 15'b100010000001011;
      12'b101101101100:
        _o_sv = 15'b100010000010000;
      12'b101101101101:
        _o_sv = 15'b100010000010101;
      12'b101101101110:
        _o_sv = 15'b100010000011011;
      12'b101101101111:
        _o_sv = 15'b100010000100000;
      12'b101101110000:
        _o_sv = 15'b100010000100101;
      12'b101101110001:
        _o_sv = 15'b100010000101011;
      12'b101101110010:
        _o_sv = 15'b100010000110000;
      12'b101101110011:
        _o_sv = 15'b100010000110101;
      12'b101101110100:
        _o_sv = 15'b100010000111011;
      12'b101101110101:
        _o_sv = 15'b100010001000000;
      12'b101101110110:
        _o_sv = 15'b100010001000101;
      12'b101101110111:
        _o_sv = 15'b100010001001011;
      12'b101101111000:
        _o_sv = 15'b100010001010000;
      12'b101101111001:
        _o_sv = 15'b100010001010101;
      12'b101101111010:
        _o_sv = 15'b100010001011010;
      12'b101101111011:
        _o_sv = 15'b100010001100000;
      12'b101101111100:
        _o_sv = 15'b100010001100101;
      12'b101101111101:
        _o_sv = 15'b100010001101010;
      12'b101101111110:
        _o_sv = 15'b100010001110000;
      12'b101101111111:
        _o_sv = 15'b100010001110101;
      12'b101110000000:
        _o_sv = 15'b100010001111010;
      12'b101110000001:
        _o_sv = 15'b100010010000000;
      12'b101110000010:
        _o_sv = 15'b100010010000101;
      12'b101110000011:
        _o_sv = 15'b100010010001010;
      12'b101110000100:
        _o_sv = 15'b100010010010000;
      12'b101110000101:
        _o_sv = 15'b100010010010101;
      12'b101110000110:
        _o_sv = 15'b100010010011010;
      12'b101110000111:
        _o_sv = 15'b100010010011111;
      12'b101110001000:
        _o_sv = 15'b100010010100101;
      12'b101110001001:
        _o_sv = 15'b100010010101010;
      12'b101110001010:
        _o_sv = 15'b100010010101111;
      12'b101110001011:
        _o_sv = 15'b100010010110101;
      12'b101110001100:
        _o_sv = 15'b100010010111010;
      12'b101110001101:
        _o_sv = 15'b100010010111111;
      12'b101110001110:
        _o_sv = 15'b100010011000101;
      12'b101110001111:
        _o_sv = 15'b100010011001010;
      12'b101110010000:
        _o_sv = 15'b100010011001111;
      12'b101110010001:
        _o_sv = 15'b100010011010100;
      12'b101110010010:
        _o_sv = 15'b100010011011010;
      12'b101110010011:
        _o_sv = 15'b100010011011111;
      12'b101110010100:
        _o_sv = 15'b100010011100100;
      12'b101110010101:
        _o_sv = 15'b100010011101010;
      12'b101110010110:
        _o_sv = 15'b100010011101111;
      12'b101110010111:
        _o_sv = 15'b100010011110100;
      12'b101110011000:
        _o_sv = 15'b100010011111010;
      12'b101110011001:
        _o_sv = 15'b100010011111111;
      12'b101110011010:
        _o_sv = 15'b100010100000100;
      12'b101110011011:
        _o_sv = 15'b100010100001001;
      12'b101110011100:
        _o_sv = 15'b100010100001111;
      12'b101110011101:
        _o_sv = 15'b100010100010100;
      12'b101110011110:
        _o_sv = 15'b100010100011001;
      12'b101110011111:
        _o_sv = 15'b100010100011111;
      12'b101110100000:
        _o_sv = 15'b100010100100100;
      12'b101110100001:
        _o_sv = 15'b100010100101001;
      12'b101110100010:
        _o_sv = 15'b100010100101110;
      12'b101110100011:
        _o_sv = 15'b100010100110100;
      12'b101110100100:
        _o_sv = 15'b100010100111001;
      12'b101110100101:
        _o_sv = 15'b100010100111110;
      12'b101110100110:
        _o_sv = 15'b100010101000100;
      12'b101110100111:
        _o_sv = 15'b100010101001001;
      12'b101110101000:
        _o_sv = 15'b100010101001110;
      12'b101110101001:
        _o_sv = 15'b100010101010011;
      12'b101110101010:
        _o_sv = 15'b100010101011001;
      12'b101110101011:
        _o_sv = 15'b100010101011110;
      12'b101110101100:
        _o_sv = 15'b100010101100011;
      12'b101110101101:
        _o_sv = 15'b100010101101001;
      12'b101110101110:
        _o_sv = 15'b100010101101110;
      12'b101110101111:
        _o_sv = 15'b100010101110011;
      12'b101110110000:
        _o_sv = 15'b100010101111000;
      12'b101110110001:
        _o_sv = 15'b100010101111110;
      12'b101110110010:
        _o_sv = 15'b100010110000011;
      12'b101110110011:
        _o_sv = 15'b100010110001000;
      12'b101110110100:
        _o_sv = 15'b100010110001101;
      12'b101110110101:
        _o_sv = 15'b100010110010011;
      12'b101110110110:
        _o_sv = 15'b100010110011000;
      12'b101110110111:
        _o_sv = 15'b100010110011101;
      12'b101110111000:
        _o_sv = 15'b100010110100011;
      12'b101110111001:
        _o_sv = 15'b100010110101000;
      12'b101110111010:
        _o_sv = 15'b100010110101101;
      12'b101110111011:
        _o_sv = 15'b100010110110010;
      12'b101110111100:
        _o_sv = 15'b100010110111000;
      12'b101110111101:
        _o_sv = 15'b100010110111101;
      12'b101110111110:
        _o_sv = 15'b100010111000010;
      12'b101110111111:
        _o_sv = 15'b100010111000111;
      12'b101111000000:
        _o_sv = 15'b100010111001101;
      12'b101111000001:
        _o_sv = 15'b100010111010010;
      12'b101111000010:
        _o_sv = 15'b100010111010111;
      12'b101111000011:
        _o_sv = 15'b100010111011101;
      12'b101111000100:
        _o_sv = 15'b100010111100010;
      12'b101111000101:
        _o_sv = 15'b100010111100111;
      12'b101111000110:
        _o_sv = 15'b100010111101100;
      12'b101111000111:
        _o_sv = 15'b100010111110010;
      12'b101111001000:
        _o_sv = 15'b100010111110111;
      12'b101111001001:
        _o_sv = 15'b100010111111100;
      12'b101111001010:
        _o_sv = 15'b100011000000001;
      12'b101111001011:
        _o_sv = 15'b100011000000111;
      12'b101111001100:
        _o_sv = 15'b100011000001100;
      12'b101111001101:
        _o_sv = 15'b100011000010001;
      12'b101111001110:
        _o_sv = 15'b100011000010110;
      12'b101111001111:
        _o_sv = 15'b100011000011100;
      12'b101111010000:
        _o_sv = 15'b100011000100001;
      12'b101111010001:
        _o_sv = 15'b100011000100110;
      12'b101111010010:
        _o_sv = 15'b100011000101011;
      12'b101111010011:
        _o_sv = 15'b100011000110001;
      12'b101111010100:
        _o_sv = 15'b100011000110110;
      12'b101111010101:
        _o_sv = 15'b100011000111011;
      12'b101111010110:
        _o_sv = 15'b100011001000000;
      12'b101111010111:
        _o_sv = 15'b100011001000110;
      12'b101111011000:
        _o_sv = 15'b100011001001011;
      12'b101111011001:
        _o_sv = 15'b100011001010000;
      12'b101111011010:
        _o_sv = 15'b100011001010101;
      12'b101111011011:
        _o_sv = 15'b100011001011011;
      12'b101111011100:
        _o_sv = 15'b100011001100000;
      12'b101111011101:
        _o_sv = 15'b100011001100101;
      12'b101111011110:
        _o_sv = 15'b100011001101010;
      12'b101111011111:
        _o_sv = 15'b100011001110000;
      12'b101111100000:
        _o_sv = 15'b100011001110101;
      12'b101111100001:
        _o_sv = 15'b100011001111010;
      12'b101111100010:
        _o_sv = 15'b100011001111111;
      12'b101111100011:
        _o_sv = 15'b100011010000101;
      12'b101111100100:
        _o_sv = 15'b100011010001010;
      12'b101111100101:
        _o_sv = 15'b100011010001111;
      12'b101111100110:
        _o_sv = 15'b100011010010100;
      12'b101111100111:
        _o_sv = 15'b100011010011010;
      12'b101111101000:
        _o_sv = 15'b100011010011111;
      12'b101111101001:
        _o_sv = 15'b100011010100100;
      12'b101111101010:
        _o_sv = 15'b100011010101001;
      12'b101111101011:
        _o_sv = 15'b100011010101111;
      12'b101111101100:
        _o_sv = 15'b100011010110100;
      12'b101111101101:
        _o_sv = 15'b100011010111001;
      12'b101111101110:
        _o_sv = 15'b100011010111110;
      12'b101111101111:
        _o_sv = 15'b100011011000100;
      12'b101111110000:
        _o_sv = 15'b100011011001001;
      12'b101111110001:
        _o_sv = 15'b100011011001110;
      12'b101111110010:
        _o_sv = 15'b100011011010011;
      12'b101111110011:
        _o_sv = 15'b100011011011000;
      12'b101111110100:
        _o_sv = 15'b100011011011110;
      12'b101111110101:
        _o_sv = 15'b100011011100011;
      12'b101111110110:
        _o_sv = 15'b100011011101000;
      12'b101111110111:
        _o_sv = 15'b100011011101101;
      12'b101111111000:
        _o_sv = 15'b100011011110011;
      12'b101111111001:
        _o_sv = 15'b100011011111000;
      12'b101111111010:
        _o_sv = 15'b100011011111101;
      12'b101111111011:
        _o_sv = 15'b100011100000010;
      12'b101111111100:
        _o_sv = 15'b100011100001000;
      12'b101111111101:
        _o_sv = 15'b100011100001101;
      12'b101111111110:
        _o_sv = 15'b100011100010010;
      12'b101111111111:
        _o_sv = 15'b100011100010111;
      12'b110000000000:
        _o_sv = 15'b100011100011100;
      12'b110000000001:
        _o_sv = 15'b100011100100010;
      12'b110000000010:
        _o_sv = 15'b100011100100111;
      12'b110000000011:
        _o_sv = 15'b100011100101100;
      12'b110000000100:
        _o_sv = 15'b100011100110001;
      12'b110000000101:
        _o_sv = 15'b100011100110111;
      12'b110000000110:
        _o_sv = 15'b100011100111100;
      12'b110000000111:
        _o_sv = 15'b100011101000001;
      12'b110000001000:
        _o_sv = 15'b100011101000110;
      12'b110000001001:
        _o_sv = 15'b100011101001011;
      12'b110000001010:
        _o_sv = 15'b100011101010001;
      12'b110000001011:
        _o_sv = 15'b100011101010110;
      12'b110000001100:
        _o_sv = 15'b100011101011011;
      12'b110000001101:
        _o_sv = 15'b100011101100000;
      12'b110000001110:
        _o_sv = 15'b100011101100101;
      12'b110000001111:
        _o_sv = 15'b100011101101011;
      12'b110000010000:
        _o_sv = 15'b100011101110000;
      12'b110000010001:
        _o_sv = 15'b100011101110101;
      12'b110000010010:
        _o_sv = 15'b100011101111010;
      12'b110000010011:
        _o_sv = 15'b100011110000000;
      12'b110000010100:
        _o_sv = 15'b100011110000101;
      12'b110000010101:
        _o_sv = 15'b100011110001010;
      12'b110000010110:
        _o_sv = 15'b100011110001111;
      12'b110000010111:
        _o_sv = 15'b100011110010100;
      12'b110000011000:
        _o_sv = 15'b100011110011010;
      12'b110000011001:
        _o_sv = 15'b100011110011111;
      12'b110000011010:
        _o_sv = 15'b100011110100100;
      12'b110000011011:
        _o_sv = 15'b100011110101001;
      12'b110000011100:
        _o_sv = 15'b100011110101110;
      12'b110000011101:
        _o_sv = 15'b100011110110100;
      12'b110000011110:
        _o_sv = 15'b100011110111001;
      12'b110000011111:
        _o_sv = 15'b100011110111110;
      12'b110000100000:
        _o_sv = 15'b100011111000011;
      12'b110000100001:
        _o_sv = 15'b100011111001000;
      12'b110000100010:
        _o_sv = 15'b100011111001110;
      12'b110000100011:
        _o_sv = 15'b100011111010011;
      12'b110000100100:
        _o_sv = 15'b100011111011000;
      12'b110000100101:
        _o_sv = 15'b100011111011101;
      12'b110000100110:
        _o_sv = 15'b100011111100010;
      12'b110000100111:
        _o_sv = 15'b100011111101000;
      12'b110000101000:
        _o_sv = 15'b100011111101101;
      12'b110000101001:
        _o_sv = 15'b100011111110010;
      12'b110000101010:
        _o_sv = 15'b100011111110111;
      12'b110000101011:
        _o_sv = 15'b100011111111100;
      12'b110000101100:
        _o_sv = 15'b100100000000010;
      12'b110000101101:
        _o_sv = 15'b100100000000111;
      12'b110000101110:
        _o_sv = 15'b100100000001100;
      12'b110000101111:
        _o_sv = 15'b100100000010001;
      12'b110000110000:
        _o_sv = 15'b100100000010110;
      12'b110000110001:
        _o_sv = 15'b100100000011100;
      12'b110000110010:
        _o_sv = 15'b100100000100001;
      12'b110000110011:
        _o_sv = 15'b100100000100110;
      12'b110000110100:
        _o_sv = 15'b100100000101011;
      12'b110000110101:
        _o_sv = 15'b100100000110000;
      12'b110000110110:
        _o_sv = 15'b100100000110110;
      12'b110000110111:
        _o_sv = 15'b100100000111011;
      12'b110000111000:
        _o_sv = 15'b100100001000000;
      12'b110000111001:
        _o_sv = 15'b100100001000101;
      12'b110000111010:
        _o_sv = 15'b100100001001010;
      12'b110000111011:
        _o_sv = 15'b100100001001111;
      12'b110000111100:
        _o_sv = 15'b100100001010101;
      12'b110000111101:
        _o_sv = 15'b100100001011010;
      12'b110000111110:
        _o_sv = 15'b100100001011111;
      12'b110000111111:
        _o_sv = 15'b100100001100100;
      12'b110001000000:
        _o_sv = 15'b100100001101001;
      12'b110001000001:
        _o_sv = 15'b100100001101111;
      12'b110001000010:
        _o_sv = 15'b100100001110100;
      12'b110001000011:
        _o_sv = 15'b100100001111001;
      12'b110001000100:
        _o_sv = 15'b100100001111110;
      12'b110001000101:
        _o_sv = 15'b100100010000011;
      12'b110001000110:
        _o_sv = 15'b100100010001000;
      12'b110001000111:
        _o_sv = 15'b100100010001110;
      12'b110001001000:
        _o_sv = 15'b100100010010011;
      12'b110001001001:
        _o_sv = 15'b100100010011000;
      12'b110001001010:
        _o_sv = 15'b100100010011101;
      12'b110001001011:
        _o_sv = 15'b100100010100010;
      12'b110001001100:
        _o_sv = 15'b100100010101000;
      12'b110001001101:
        _o_sv = 15'b100100010101101;
      12'b110001001110:
        _o_sv = 15'b100100010110010;
      12'b110001001111:
        _o_sv = 15'b100100010110111;
      12'b110001010000:
        _o_sv = 15'b100100010111100;
      12'b110001010001:
        _o_sv = 15'b100100011000001;
      12'b110001010010:
        _o_sv = 15'b100100011000111;
      12'b110001010011:
        _o_sv = 15'b100100011001100;
      12'b110001010100:
        _o_sv = 15'b100100011010001;
      12'b110001010101:
        _o_sv = 15'b100100011010110;
      12'b110001010110:
        _o_sv = 15'b100100011011011;
      12'b110001010111:
        _o_sv = 15'b100100011100000;
      12'b110001011000:
        _o_sv = 15'b100100011100110;
      12'b110001011001:
        _o_sv = 15'b100100011101011;
      12'b110001011010:
        _o_sv = 15'b100100011110000;
      12'b110001011011:
        _o_sv = 15'b100100011110101;
      12'b110001011100:
        _o_sv = 15'b100100011111010;
      12'b110001011101:
        _o_sv = 15'b100100011111111;
      12'b110001011110:
        _o_sv = 15'b100100100000101;
      12'b110001011111:
        _o_sv = 15'b100100100001010;
      12'b110001100000:
        _o_sv = 15'b100100100001111;
      12'b110001100001:
        _o_sv = 15'b100100100010100;
      12'b110001100010:
        _o_sv = 15'b100100100011001;
      12'b110001100011:
        _o_sv = 15'b100100100011110;
      12'b110001100100:
        _o_sv = 15'b100100100100011;
      12'b110001100101:
        _o_sv = 15'b100100100101001;
      12'b110001100110:
        _o_sv = 15'b100100100101110;
      12'b110001100111:
        _o_sv = 15'b100100100110011;
      12'b110001101000:
        _o_sv = 15'b100100100111000;
      12'b110001101001:
        _o_sv = 15'b100100100111101;
      12'b110001101010:
        _o_sv = 15'b100100101000010;
      12'b110001101011:
        _o_sv = 15'b100100101001000;
      12'b110001101100:
        _o_sv = 15'b100100101001101;
      12'b110001101101:
        _o_sv = 15'b100100101010010;
      12'b110001101110:
        _o_sv = 15'b100100101010111;
      12'b110001101111:
        _o_sv = 15'b100100101011100;
      12'b110001110000:
        _o_sv = 15'b100100101100001;
      12'b110001110001:
        _o_sv = 15'b100100101100110;
      12'b110001110010:
        _o_sv = 15'b100100101101100;
      12'b110001110011:
        _o_sv = 15'b100100101110001;
      12'b110001110100:
        _o_sv = 15'b100100101110110;
      12'b110001110101:
        _o_sv = 15'b100100101111011;
      12'b110001110110:
        _o_sv = 15'b100100110000000;
      12'b110001110111:
        _o_sv = 15'b100100110000101;
      12'b110001111000:
        _o_sv = 15'b100100110001010;
      12'b110001111001:
        _o_sv = 15'b100100110010000;
      12'b110001111010:
        _o_sv = 15'b100100110010101;
      12'b110001111011:
        _o_sv = 15'b100100110011010;
      12'b110001111100:
        _o_sv = 15'b100100110011111;
      12'b110001111101:
        _o_sv = 15'b100100110100100;
      12'b110001111110:
        _o_sv = 15'b100100110101001;
      12'b110001111111:
        _o_sv = 15'b100100110101110;
      12'b110010000000:
        _o_sv = 15'b100100110110100;
      12'b110010000001:
        _o_sv = 15'b100100110111001;
      12'b110010000010:
        _o_sv = 15'b100100110111110;
      12'b110010000011:
        _o_sv = 15'b100100111000011;
      12'b110010000100:
        _o_sv = 15'b100100111001000;
      12'b110010000101:
        _o_sv = 15'b100100111001101;
      12'b110010000110:
        _o_sv = 15'b100100111010010;
      12'b110010000111:
        _o_sv = 15'b100100111011000;
      12'b110010001000:
        _o_sv = 15'b100100111011101;
      12'b110010001001:
        _o_sv = 15'b100100111100010;
      12'b110010001010:
        _o_sv = 15'b100100111100111;
      12'b110010001011:
        _o_sv = 15'b100100111101100;
      12'b110010001100:
        _o_sv = 15'b100100111110001;
      12'b110010001101:
        _o_sv = 15'b100100111110110;
      12'b110010001110:
        _o_sv = 15'b100100111111011;
      12'b110010001111:
        _o_sv = 15'b100101000000001;
      12'b110010010000:
        _o_sv = 15'b100101000000110;
      12'b110010010001:
        _o_sv = 15'b100101000001011;
      12'b110010010010:
        _o_sv = 15'b100101000010000;
      12'b110010010011:
        _o_sv = 15'b100101000010101;
      12'b110010010100:
        _o_sv = 15'b100101000011010;
      12'b110010010101:
        _o_sv = 15'b100101000011111;
      12'b110010010110:
        _o_sv = 15'b100101000100100;
      12'b110010010111:
        _o_sv = 15'b100101000101010;
      12'b110010011000:
        _o_sv = 15'b100101000101111;
      12'b110010011001:
        _o_sv = 15'b100101000110100;
      12'b110010011010:
        _o_sv = 15'b100101000111001;
      12'b110010011011:
        _o_sv = 15'b100101000111110;
      12'b110010011100:
        _o_sv = 15'b100101001000011;
      12'b110010011101:
        _o_sv = 15'b100101001001000;
      12'b110010011110:
        _o_sv = 15'b100101001001101;
      12'b110010011111:
        _o_sv = 15'b100101001010010;
      12'b110010100000:
        _o_sv = 15'b100101001011000;
      12'b110010100001:
        _o_sv = 15'b100101001011101;
      12'b110010100010:
        _o_sv = 15'b100101001100010;
      12'b110010100011:
        _o_sv = 15'b100101001100111;
      12'b110010100100:
        _o_sv = 15'b100101001101100;
      12'b110010100101:
        _o_sv = 15'b100101001110001;
      12'b110010100110:
        _o_sv = 15'b100101001110110;
      12'b110010100111:
        _o_sv = 15'b100101001111011;
      12'b110010101000:
        _o_sv = 15'b100101010000001;
      12'b110010101001:
        _o_sv = 15'b100101010000110;
      12'b110010101010:
        _o_sv = 15'b100101010001011;
      12'b110010101011:
        _o_sv = 15'b100101010010000;
      12'b110010101100:
        _o_sv = 15'b100101010010101;
      12'b110010101101:
        _o_sv = 15'b100101010011010;
      12'b110010101110:
        _o_sv = 15'b100101010011111;
      12'b110010101111:
        _o_sv = 15'b100101010100100;
      12'b110010110000:
        _o_sv = 15'b100101010101001;
      12'b110010110001:
        _o_sv = 15'b100101010101110;
      12'b110010110010:
        _o_sv = 15'b100101010110100;
      12'b110010110011:
        _o_sv = 15'b100101010111001;
      12'b110010110100:
        _o_sv = 15'b100101010111110;
      12'b110010110101:
        _o_sv = 15'b100101011000011;
      12'b110010110110:
        _o_sv = 15'b100101011001000;
      12'b110010110111:
        _o_sv = 15'b100101011001101;
      12'b110010111000:
        _o_sv = 15'b100101011010010;
      12'b110010111001:
        _o_sv = 15'b100101011010111;
      12'b110010111010:
        _o_sv = 15'b100101011011100;
      12'b110010111011:
        _o_sv = 15'b100101011100001;
      12'b110010111100:
        _o_sv = 15'b100101011100111;
      12'b110010111101:
        _o_sv = 15'b100101011101100;
      12'b110010111110:
        _o_sv = 15'b100101011110001;
      12'b110010111111:
        _o_sv = 15'b100101011110110;
      12'b110011000000:
        _o_sv = 15'b100101011111011;
      12'b110011000001:
        _o_sv = 15'b100101100000000;
      12'b110011000010:
        _o_sv = 15'b100101100000101;
      12'b110011000011:
        _o_sv = 15'b100101100001010;
      12'b110011000100:
        _o_sv = 15'b100101100001111;
      12'b110011000101:
        _o_sv = 15'b100101100010100;
      12'b110011000110:
        _o_sv = 15'b100101100011001;
      12'b110011000111:
        _o_sv = 15'b100101100011111;
      12'b110011001000:
        _o_sv = 15'b100101100100100;
      12'b110011001001:
        _o_sv = 15'b100101100101001;
      12'b110011001010:
        _o_sv = 15'b100101100101110;
      12'b110011001011:
        _o_sv = 15'b100101100110011;
      12'b110011001100:
        _o_sv = 15'b100101100111000;
      12'b110011001101:
        _o_sv = 15'b100101100111101;
      12'b110011001110:
        _o_sv = 15'b100101101000010;
      12'b110011001111:
        _o_sv = 15'b100101101000111;
      12'b110011010000:
        _o_sv = 15'b100101101001100;
      12'b110011010001:
        _o_sv = 15'b100101101010001;
      12'b110011010010:
        _o_sv = 15'b100101101010110;
      12'b110011010011:
        _o_sv = 15'b100101101011100;
      12'b110011010100:
        _o_sv = 15'b100101101100001;
      12'b110011010101:
        _o_sv = 15'b100101101100110;
      12'b110011010110:
        _o_sv = 15'b100101101101011;
      12'b110011010111:
        _o_sv = 15'b100101101110000;
      12'b110011011000:
        _o_sv = 15'b100101101110101;
      12'b110011011001:
        _o_sv = 15'b100101101111010;
      12'b110011011010:
        _o_sv = 15'b100101101111111;
      12'b110011011011:
        _o_sv = 15'b100101110000100;
      12'b110011011100:
        _o_sv = 15'b100101110001001;
      12'b110011011101:
        _o_sv = 15'b100101110001110;
      12'b110011011110:
        _o_sv = 15'b100101110010011;
      12'b110011011111:
        _o_sv = 15'b100101110011000;
      12'b110011100000:
        _o_sv = 15'b100101110011110;
      12'b110011100001:
        _o_sv = 15'b100101110100011;
      12'b110011100010:
        _o_sv = 15'b100101110101000;
      12'b110011100011:
        _o_sv = 15'b100101110101101;
      12'b110011100100:
        _o_sv = 15'b100101110110010;
      12'b110011100101:
        _o_sv = 15'b100101110110111;
      12'b110011100110:
        _o_sv = 15'b100101110111100;
      12'b110011100111:
        _o_sv = 15'b100101111000001;
      12'b110011101000:
        _o_sv = 15'b100101111000110;
      12'b110011101001:
        _o_sv = 15'b100101111001011;
      12'b110011101010:
        _o_sv = 15'b100101111010000;
      12'b110011101011:
        _o_sv = 15'b100101111010101;
      12'b110011101100:
        _o_sv = 15'b100101111011010;
      12'b110011101101:
        _o_sv = 15'b100101111011111;
      12'b110011101110:
        _o_sv = 15'b100101111100100;
      12'b110011101111:
        _o_sv = 15'b100101111101001;
      12'b110011110000:
        _o_sv = 15'b100101111101111;
      12'b110011110001:
        _o_sv = 15'b100101111110100;
      12'b110011110010:
        _o_sv = 15'b100101111111001;
      12'b110011110011:
        _o_sv = 15'b100101111111110;
      12'b110011110100:
        _o_sv = 15'b100110000000011;
      12'b110011110101:
        _o_sv = 15'b100110000001000;
      12'b110011110110:
        _o_sv = 15'b100110000001101;
      12'b110011110111:
        _o_sv = 15'b100110000010010;
      12'b110011111000:
        _o_sv = 15'b100110000010111;
      12'b110011111001:
        _o_sv = 15'b100110000011100;
      12'b110011111010:
        _o_sv = 15'b100110000100001;
      12'b110011111011:
        _o_sv = 15'b100110000100110;
      12'b110011111100:
        _o_sv = 15'b100110000101011;
      12'b110011111101:
        _o_sv = 15'b100110000110000;
      12'b110011111110:
        _o_sv = 15'b100110000110101;
      12'b110011111111:
        _o_sv = 15'b100110000111010;
      12'b110100000000:
        _o_sv = 15'b100110000111111;
      12'b110100000001:
        _o_sv = 15'b100110001000100;
      12'b110100000010:
        _o_sv = 15'b100110001001001;
      12'b110100000011:
        _o_sv = 15'b100110001001111;
      12'b110100000100:
        _o_sv = 15'b100110001010100;
      12'b110100000101:
        _o_sv = 15'b100110001011001;
      12'b110100000110:
        _o_sv = 15'b100110001011110;
      12'b110100000111:
        _o_sv = 15'b100110001100011;
      12'b110100001000:
        _o_sv = 15'b100110001101000;
      12'b110100001001:
        _o_sv = 15'b100110001101101;
      12'b110100001010:
        _o_sv = 15'b100110001110010;
      12'b110100001011:
        _o_sv = 15'b100110001110111;
      12'b110100001100:
        _o_sv = 15'b100110001111100;
      12'b110100001101:
        _o_sv = 15'b100110010000001;
      12'b110100001110:
        _o_sv = 15'b100110010000110;
      12'b110100001111:
        _o_sv = 15'b100110010001011;
      12'b110100010000:
        _o_sv = 15'b100110010010000;
      12'b110100010001:
        _o_sv = 15'b100110010010101;
      12'b110100010010:
        _o_sv = 15'b100110010011010;
      12'b110100010011:
        _o_sv = 15'b100110010011111;
      12'b110100010100:
        _o_sv = 15'b100110010100100;
      12'b110100010101:
        _o_sv = 15'b100110010101001;
      12'b110100010110:
        _o_sv = 15'b100110010101110;
      12'b110100010111:
        _o_sv = 15'b100110010110011;
      12'b110100011000:
        _o_sv = 15'b100110010111000;
      12'b110100011001:
        _o_sv = 15'b100110010111101;
      12'b110100011010:
        _o_sv = 15'b100110011000010;
      12'b110100011011:
        _o_sv = 15'b100110011000111;
      12'b110100011100:
        _o_sv = 15'b100110011001100;
      12'b110100011101:
        _o_sv = 15'b100110011010001;
      12'b110100011110:
        _o_sv = 15'b100110011010110;
      12'b110100011111:
        _o_sv = 15'b100110011011011;
      12'b110100100000:
        _o_sv = 15'b100110011100001;
      12'b110100100001:
        _o_sv = 15'b100110011100110;
      12'b110100100010:
        _o_sv = 15'b100110011101011;
      12'b110100100011:
        _o_sv = 15'b100110011110000;
      12'b110100100100:
        _o_sv = 15'b100110011110101;
      12'b110100100101:
        _o_sv = 15'b100110011111010;
      12'b110100100110:
        _o_sv = 15'b100110011111111;
      12'b110100100111:
        _o_sv = 15'b100110100000100;
      12'b110100101000:
        _o_sv = 15'b100110100001001;
      12'b110100101001:
        _o_sv = 15'b100110100001110;
      12'b110100101010:
        _o_sv = 15'b100110100010011;
      12'b110100101011:
        _o_sv = 15'b100110100011000;
      12'b110100101100:
        _o_sv = 15'b100110100011101;
      12'b110100101101:
        _o_sv = 15'b100110100100010;
      12'b110100101110:
        _o_sv = 15'b100110100100111;
      12'b110100101111:
        _o_sv = 15'b100110100101100;
      12'b110100110000:
        _o_sv = 15'b100110100110001;
      12'b110100110001:
        _o_sv = 15'b100110100110110;
      12'b110100110010:
        _o_sv = 15'b100110100111011;
      12'b110100110011:
        _o_sv = 15'b100110101000000;
      12'b110100110100:
        _o_sv = 15'b100110101000101;
      12'b110100110101:
        _o_sv = 15'b100110101001010;
      12'b110100110110:
        _o_sv = 15'b100110101001111;
      12'b110100110111:
        _o_sv = 15'b100110101010100;
      12'b110100111000:
        _o_sv = 15'b100110101011001;
      12'b110100111001:
        _o_sv = 15'b100110101011110;
      12'b110100111010:
        _o_sv = 15'b100110101100011;
      12'b110100111011:
        _o_sv = 15'b100110101101000;
      12'b110100111100:
        _o_sv = 15'b100110101101101;
      12'b110100111101:
        _o_sv = 15'b100110101110010;
      12'b110100111110:
        _o_sv = 15'b100110101110111;
      12'b110100111111:
        _o_sv = 15'b100110101111100;
      12'b110101000000:
        _o_sv = 15'b100110110000001;
      12'b110101000001:
        _o_sv = 15'b100110110000110;
      12'b110101000010:
        _o_sv = 15'b100110110001011;
      12'b110101000011:
        _o_sv = 15'b100110110010000;
      12'b110101000100:
        _o_sv = 15'b100110110010101;
      12'b110101000101:
        _o_sv = 15'b100110110011010;
      12'b110101000110:
        _o_sv = 15'b100110110011111;
      12'b110101000111:
        _o_sv = 15'b100110110100100;
      12'b110101001000:
        _o_sv = 15'b100110110101001;
      12'b110101001001:
        _o_sv = 15'b100110110101110;
      12'b110101001010:
        _o_sv = 15'b100110110110011;
      12'b110101001011:
        _o_sv = 15'b100110110111000;
      12'b110101001100:
        _o_sv = 15'b100110110111101;
      12'b110101001101:
        _o_sv = 15'b100110111000010;
      12'b110101001110:
        _o_sv = 15'b100110111000111;
      12'b110101001111:
        _o_sv = 15'b100110111001100;
      12'b110101010000:
        _o_sv = 15'b100110111010001;
      12'b110101010001:
        _o_sv = 15'b100110111010110;
      12'b110101010010:
        _o_sv = 15'b100110111011011;
      12'b110101010011:
        _o_sv = 15'b100110111100000;
      12'b110101010100:
        _o_sv = 15'b100110111100101;
      12'b110101010101:
        _o_sv = 15'b100110111101010;
      12'b110101010110:
        _o_sv = 15'b100110111101111;
      12'b110101010111:
        _o_sv = 15'b100110111110100;
      12'b110101011000:
        _o_sv = 15'b100110111111001;
      12'b110101011001:
        _o_sv = 15'b100110111111110;
      12'b110101011010:
        _o_sv = 15'b100111000000011;
      12'b110101011011:
        _o_sv = 15'b100111000001000;
      12'b110101011100:
        _o_sv = 15'b100111000001101;
      12'b110101011101:
        _o_sv = 15'b100111000010010;
      12'b110101011110:
        _o_sv = 15'b100111000010111;
      12'b110101011111:
        _o_sv = 15'b100111000011100;
      12'b110101100000:
        _o_sv = 15'b100111000100001;
      12'b110101100001:
        _o_sv = 15'b100111000100110;
      12'b110101100010:
        _o_sv = 15'b100111000101010;
      12'b110101100011:
        _o_sv = 15'b100111000101111;
      12'b110101100100:
        _o_sv = 15'b100111000110100;
      12'b110101100101:
        _o_sv = 15'b100111000111001;
      12'b110101100110:
        _o_sv = 15'b100111000111110;
      12'b110101100111:
        _o_sv = 15'b100111001000011;
      12'b110101101000:
        _o_sv = 15'b100111001001000;
      12'b110101101001:
        _o_sv = 15'b100111001001101;
      12'b110101101010:
        _o_sv = 15'b100111001010010;
      12'b110101101011:
        _o_sv = 15'b100111001010111;
      12'b110101101100:
        _o_sv = 15'b100111001011100;
      12'b110101101101:
        _o_sv = 15'b100111001100001;
      12'b110101101110:
        _o_sv = 15'b100111001100110;
      12'b110101101111:
        _o_sv = 15'b100111001101011;
      12'b110101110000:
        _o_sv = 15'b100111001110000;
      12'b110101110001:
        _o_sv = 15'b100111001110101;
      12'b110101110010:
        _o_sv = 15'b100111001111010;
      12'b110101110011:
        _o_sv = 15'b100111001111111;
      12'b110101110100:
        _o_sv = 15'b100111010000100;
      12'b110101110101:
        _o_sv = 15'b100111010001001;
      12'b110101110110:
        _o_sv = 15'b100111010001110;
      12'b110101110111:
        _o_sv = 15'b100111010010011;
      12'b110101111000:
        _o_sv = 15'b100111010011000;
      12'b110101111001:
        _o_sv = 15'b100111010011101;
      12'b110101111010:
        _o_sv = 15'b100111010100010;
      12'b110101111011:
        _o_sv = 15'b100111010100111;
      12'b110101111100:
        _o_sv = 15'b100111010101100;
      12'b110101111101:
        _o_sv = 15'b100111010110001;
      12'b110101111110:
        _o_sv = 15'b100111010110110;
      12'b110101111111:
        _o_sv = 15'b100111010111010;
      12'b110110000000:
        _o_sv = 15'b100111010111111;
      12'b110110000001:
        _o_sv = 15'b100111011000100;
      12'b110110000010:
        _o_sv = 15'b100111011001001;
      12'b110110000011:
        _o_sv = 15'b100111011001110;
      12'b110110000100:
        _o_sv = 15'b100111011010011;
      12'b110110000101:
        _o_sv = 15'b100111011011000;
      12'b110110000110:
        _o_sv = 15'b100111011011101;
      12'b110110000111:
        _o_sv = 15'b100111011100010;
      12'b110110001000:
        _o_sv = 15'b100111011100111;
      12'b110110001001:
        _o_sv = 15'b100111011101100;
      12'b110110001010:
        _o_sv = 15'b100111011110001;
      12'b110110001011:
        _o_sv = 15'b100111011110110;
      12'b110110001100:
        _o_sv = 15'b100111011111011;
      12'b110110001101:
        _o_sv = 15'b100111100000000;
      12'b110110001110:
        _o_sv = 15'b100111100000101;
      12'b110110001111:
        _o_sv = 15'b100111100001010;
      12'b110110010000:
        _o_sv = 15'b100111100001111;
      12'b110110010001:
        _o_sv = 15'b100111100010100;
      12'b110110010010:
        _o_sv = 15'b100111100011000;
      12'b110110010011:
        _o_sv = 15'b100111100011101;
      12'b110110010100:
        _o_sv = 15'b100111100100010;
      12'b110110010101:
        _o_sv = 15'b100111100100111;
      12'b110110010110:
        _o_sv = 15'b100111100101100;
      12'b110110010111:
        _o_sv = 15'b100111100110001;
      12'b110110011000:
        _o_sv = 15'b100111100110110;
      12'b110110011001:
        _o_sv = 15'b100111100111011;
      12'b110110011010:
        _o_sv = 15'b100111101000000;
      12'b110110011011:
        _o_sv = 15'b100111101000101;
      12'b110110011100:
        _o_sv = 15'b100111101001010;
      12'b110110011101:
        _o_sv = 15'b100111101001111;
      12'b110110011110:
        _o_sv = 15'b100111101010100;
      12'b110110011111:
        _o_sv = 15'b100111101011001;
      12'b110110100000:
        _o_sv = 15'b100111101011110;
      12'b110110100001:
        _o_sv = 15'b100111101100010;
      12'b110110100010:
        _o_sv = 15'b100111101100111;
      12'b110110100011:
        _o_sv = 15'b100111101101100;
      12'b110110100100:
        _o_sv = 15'b100111101110001;
      12'b110110100101:
        _o_sv = 15'b100111101110110;
      12'b110110100110:
        _o_sv = 15'b100111101111011;
      12'b110110100111:
        _o_sv = 15'b100111110000000;
      12'b110110101000:
        _o_sv = 15'b100111110000101;
      12'b110110101001:
        _o_sv = 15'b100111110001010;
      12'b110110101010:
        _o_sv = 15'b100111110001111;
      12'b110110101011:
        _o_sv = 15'b100111110010100;
      12'b110110101100:
        _o_sv = 15'b100111110011001;
      12'b110110101101:
        _o_sv = 15'b100111110011110;
      12'b110110101110:
        _o_sv = 15'b100111110100010;
      12'b110110101111:
        _o_sv = 15'b100111110100111;
      12'b110110110000:
        _o_sv = 15'b100111110101100;
      12'b110110110001:
        _o_sv = 15'b100111110110001;
      12'b110110110010:
        _o_sv = 15'b100111110110110;
      12'b110110110011:
        _o_sv = 15'b100111110111011;
      12'b110110110100:
        _o_sv = 15'b100111111000000;
      12'b110110110101:
        _o_sv = 15'b100111111000101;
      12'b110110110110:
        _o_sv = 15'b100111111001010;
      12'b110110110111:
        _o_sv = 15'b100111111001111;
      12'b110110111000:
        _o_sv = 15'b100111111010100;
      12'b110110111001:
        _o_sv = 15'b100111111011001;
      12'b110110111010:
        _o_sv = 15'b100111111011101;
      12'b110110111011:
        _o_sv = 15'b100111111100010;
      12'b110110111100:
        _o_sv = 15'b100111111100111;
      12'b110110111101:
        _o_sv = 15'b100111111101100;
      12'b110110111110:
        _o_sv = 15'b100111111110001;
      12'b110110111111:
        _o_sv = 15'b100111111110110;
      12'b110111000000:
        _o_sv = 15'b100111111111011;
      12'b110111000001:
        _o_sv = 15'b101000000000000;
      12'b110111000010:
        _o_sv = 15'b101000000000101;
      12'b110111000011:
        _o_sv = 15'b101000000001010;
      12'b110111000100:
        _o_sv = 15'b101000000001111;
      12'b110111000101:
        _o_sv = 15'b101000000010011;
      12'b110111000110:
        _o_sv = 15'b101000000011000;
      12'b110111000111:
        _o_sv = 15'b101000000011101;
      12'b110111001000:
        _o_sv = 15'b101000000100010;
      12'b110111001001:
        _o_sv = 15'b101000000100111;
      12'b110111001010:
        _o_sv = 15'b101000000101100;
      12'b110111001011:
        _o_sv = 15'b101000000110001;
      12'b110111001100:
        _o_sv = 15'b101000000110110;
      12'b110111001101:
        _o_sv = 15'b101000000111011;
      12'b110111001110:
        _o_sv = 15'b101000000111111;
      12'b110111001111:
        _o_sv = 15'b101000001000100;
      12'b110111010000:
        _o_sv = 15'b101000001001001;
      12'b110111010001:
        _o_sv = 15'b101000001001110;
      12'b110111010010:
        _o_sv = 15'b101000001010011;
      12'b110111010011:
        _o_sv = 15'b101000001011000;
      12'b110111010100:
        _o_sv = 15'b101000001011101;
      12'b110111010101:
        _o_sv = 15'b101000001100010;
      12'b110111010110:
        _o_sv = 15'b101000001100111;
      12'b110111010111:
        _o_sv = 15'b101000001101100;
      12'b110111011000:
        _o_sv = 15'b101000001110000;
      12'b110111011001:
        _o_sv = 15'b101000001110101;
      12'b110111011010:
        _o_sv = 15'b101000001111010;
      12'b110111011011:
        _o_sv = 15'b101000001111111;
      12'b110111011100:
        _o_sv = 15'b101000010000100;
      12'b110111011101:
        _o_sv = 15'b101000010001001;
      12'b110111011110:
        _o_sv = 15'b101000010001110;
      12'b110111011111:
        _o_sv = 15'b101000010010011;
      12'b110111100000:
        _o_sv = 15'b101000010010111;
      12'b110111100001:
        _o_sv = 15'b101000010011100;
      12'b110111100010:
        _o_sv = 15'b101000010100001;
      12'b110111100011:
        _o_sv = 15'b101000010100110;
      12'b110111100100:
        _o_sv = 15'b101000010101011;
      12'b110111100101:
        _o_sv = 15'b101000010110000;
      12'b110111100110:
        _o_sv = 15'b101000010110101;
      12'b110111100111:
        _o_sv = 15'b101000010111010;
      12'b110111101000:
        _o_sv = 15'b101000010111111;
      12'b110111101001:
        _o_sv = 15'b101000011000011;
      12'b110111101010:
        _o_sv = 15'b101000011001000;
      12'b110111101011:
        _o_sv = 15'b101000011001101;
      12'b110111101100:
        _o_sv = 15'b101000011010010;
      12'b110111101101:
        _o_sv = 15'b101000011010111;
      12'b110111101110:
        _o_sv = 15'b101000011011100;
      12'b110111101111:
        _o_sv = 15'b101000011100001;
      12'b110111110000:
        _o_sv = 15'b101000011100101;
      12'b110111110001:
        _o_sv = 15'b101000011101010;
      12'b110111110010:
        _o_sv = 15'b101000011101111;
      12'b110111110011:
        _o_sv = 15'b101000011110100;
      12'b110111110100:
        _o_sv = 15'b101000011111001;
      12'b110111110101:
        _o_sv = 15'b101000011111110;
      12'b110111110110:
        _o_sv = 15'b101000100000011;
      12'b110111110111:
        _o_sv = 15'b101000100001000;
      12'b110111111000:
        _o_sv = 15'b101000100001100;
      12'b110111111001:
        _o_sv = 15'b101000100010001;
      12'b110111111010:
        _o_sv = 15'b101000100010110;
      12'b110111111011:
        _o_sv = 15'b101000100011011;
      12'b110111111100:
        _o_sv = 15'b101000100100000;
      12'b110111111101:
        _o_sv = 15'b101000100100101;
      12'b110111111110:
        _o_sv = 15'b101000100101010;
      12'b110111111111:
        _o_sv = 15'b101000100101110;
      12'b111000000000:
        _o_sv = 15'b101000100110011;
      12'b111000000001:
        _o_sv = 15'b101000100111000;
      12'b111000000010:
        _o_sv = 15'b101000100111101;
      12'b111000000011:
        _o_sv = 15'b101000101000010;
      12'b111000000100:
        _o_sv = 15'b101000101000111;
      12'b111000000101:
        _o_sv = 15'b101000101001100;
      12'b111000000110:
        _o_sv = 15'b101000101010000;
      12'b111000000111:
        _o_sv = 15'b101000101010101;
      12'b111000001000:
        _o_sv = 15'b101000101011010;
      12'b111000001001:
        _o_sv = 15'b101000101011111;
      12'b111000001010:
        _o_sv = 15'b101000101100100;
      12'b111000001011:
        _o_sv = 15'b101000101101001;
      12'b111000001100:
        _o_sv = 15'b101000101101110;
      12'b111000001101:
        _o_sv = 15'b101000101110010;
      12'b111000001110:
        _o_sv = 15'b101000101110111;
      12'b111000001111:
        _o_sv = 15'b101000101111100;
      12'b111000010000:
        _o_sv = 15'b101000110000001;
      12'b111000010001:
        _o_sv = 15'b101000110000110;
      12'b111000010010:
        _o_sv = 15'b101000110001011;
      12'b111000010011:
        _o_sv = 15'b101000110001111;
      12'b111000010100:
        _o_sv = 15'b101000110010100;
      12'b111000010101:
        _o_sv = 15'b101000110011001;
      12'b111000010110:
        _o_sv = 15'b101000110011110;
      12'b111000010111:
        _o_sv = 15'b101000110100011;
      12'b111000011000:
        _o_sv = 15'b101000110101000;
      12'b111000011001:
        _o_sv = 15'b101000110101100;
      12'b111000011010:
        _o_sv = 15'b101000110110001;
      12'b111000011011:
        _o_sv = 15'b101000110110110;
      12'b111000011100:
        _o_sv = 15'b101000110111011;
      12'b111000011101:
        _o_sv = 15'b101000111000000;
      12'b111000011110:
        _o_sv = 15'b101000111000101;
      12'b111000011111:
        _o_sv = 15'b101000111001001;
      12'b111000100000:
        _o_sv = 15'b101000111001110;
      12'b111000100001:
        _o_sv = 15'b101000111010011;
      12'b111000100010:
        _o_sv = 15'b101000111011000;
      12'b111000100011:
        _o_sv = 15'b101000111011101;
      12'b111000100100:
        _o_sv = 15'b101000111100010;
      12'b111000100101:
        _o_sv = 15'b101000111100110;
      12'b111000100110:
        _o_sv = 15'b101000111101011;
      12'b111000100111:
        _o_sv = 15'b101000111110000;
      12'b111000101000:
        _o_sv = 15'b101000111110101;
      12'b111000101001:
        _o_sv = 15'b101000111111010;
      12'b111000101010:
        _o_sv = 15'b101000111111111;
      12'b111000101011:
        _o_sv = 15'b101001000000011;
      12'b111000101100:
        _o_sv = 15'b101001000001000;
      12'b111000101101:
        _o_sv = 15'b101001000001101;
      12'b111000101110:
        _o_sv = 15'b101001000010010;
      12'b111000101111:
        _o_sv = 15'b101001000010111;
      12'b111000110000:
        _o_sv = 15'b101001000011100;
      12'b111000110001:
        _o_sv = 15'b101001000100000;
      12'b111000110010:
        _o_sv = 15'b101001000100101;
      12'b111000110011:
        _o_sv = 15'b101001000101010;
      12'b111000110100:
        _o_sv = 15'b101001000101111;
      12'b111000110101:
        _o_sv = 15'b101001000110100;
      12'b111000110110:
        _o_sv = 15'b101001000111000;
      12'b111000110111:
        _o_sv = 15'b101001000111101;
      12'b111000111000:
        _o_sv = 15'b101001001000010;
      12'b111000111001:
        _o_sv = 15'b101001001000111;
      12'b111000111010:
        _o_sv = 15'b101001001001100;
      12'b111000111011:
        _o_sv = 15'b101001001010001;
      12'b111000111100:
        _o_sv = 15'b101001001010101;
      12'b111000111101:
        _o_sv = 15'b101001001011010;
      12'b111000111110:
        _o_sv = 15'b101001001011111;
      12'b111000111111:
        _o_sv = 15'b101001001100100;
      12'b111001000000:
        _o_sv = 15'b101001001101001;
      12'b111001000001:
        _o_sv = 15'b101001001101101;
      12'b111001000010:
        _o_sv = 15'b101001001110010;
      12'b111001000011:
        _o_sv = 15'b101001001110111;
      12'b111001000100:
        _o_sv = 15'b101001001111100;
      12'b111001000101:
        _o_sv = 15'b101001010000001;
      12'b111001000110:
        _o_sv = 15'b101001010000101;
      12'b111001000111:
        _o_sv = 15'b101001010001010;
      12'b111001001000:
        _o_sv = 15'b101001010001111;
      12'b111001001001:
        _o_sv = 15'b101001010010100;
      12'b111001001010:
        _o_sv = 15'b101001010011001;
      12'b111001001011:
        _o_sv = 15'b101001010011101;
      12'b111001001100:
        _o_sv = 15'b101001010100010;
      12'b111001001101:
        _o_sv = 15'b101001010100111;
      12'b111001001110:
        _o_sv = 15'b101001010101100;
      12'b111001001111:
        _o_sv = 15'b101001010110001;
      12'b111001010000:
        _o_sv = 15'b101001010110101;
      12'b111001010001:
        _o_sv = 15'b101001010111010;
      12'b111001010010:
        _o_sv = 15'b101001010111111;
      12'b111001010011:
        _o_sv = 15'b101001011000100;
      12'b111001010100:
        _o_sv = 15'b101001011001001;
      12'b111001010101:
        _o_sv = 15'b101001011001101;
      12'b111001010110:
        _o_sv = 15'b101001011010010;
      12'b111001010111:
        _o_sv = 15'b101001011010111;
      12'b111001011000:
        _o_sv = 15'b101001011011100;
      12'b111001011001:
        _o_sv = 15'b101001011100001;
      12'b111001011010:
        _o_sv = 15'b101001011100101;
      12'b111001011011:
        _o_sv = 15'b101001011101010;
      12'b111001011100:
        _o_sv = 15'b101001011101111;
      12'b111001011101:
        _o_sv = 15'b101001011110100;
      12'b111001011110:
        _o_sv = 15'b101001011111000;
      12'b111001011111:
        _o_sv = 15'b101001011111101;
      12'b111001100000:
        _o_sv = 15'b101001100000010;
      12'b111001100001:
        _o_sv = 15'b101001100000111;
      12'b111001100010:
        _o_sv = 15'b101001100001100;
      12'b111001100011:
        _o_sv = 15'b101001100010000;
      12'b111001100100:
        _o_sv = 15'b101001100010101;
      12'b111001100101:
        _o_sv = 15'b101001100011010;
      12'b111001100110:
        _o_sv = 15'b101001100011111;
      12'b111001100111:
        _o_sv = 15'b101001100100011;
      12'b111001101000:
        _o_sv = 15'b101001100101000;
      12'b111001101001:
        _o_sv = 15'b101001100101101;
      12'b111001101010:
        _o_sv = 15'b101001100110010;
      12'b111001101011:
        _o_sv = 15'b101001100110111;
      12'b111001101100:
        _o_sv = 15'b101001100111011;
      12'b111001101101:
        _o_sv = 15'b101001101000000;
      12'b111001101110:
        _o_sv = 15'b101001101000101;
      12'b111001101111:
        _o_sv = 15'b101001101001010;
      12'b111001110000:
        _o_sv = 15'b101001101001110;
      12'b111001110001:
        _o_sv = 15'b101001101010011;
      12'b111001110010:
        _o_sv = 15'b101001101011000;
      12'b111001110011:
        _o_sv = 15'b101001101011101;
      12'b111001110100:
        _o_sv = 15'b101001101100010;
      12'b111001110101:
        _o_sv = 15'b101001101100110;
      12'b111001110110:
        _o_sv = 15'b101001101101011;
      12'b111001110111:
        _o_sv = 15'b101001101110000;
      12'b111001111000:
        _o_sv = 15'b101001101110101;
      12'b111001111001:
        _o_sv = 15'b101001101111001;
      12'b111001111010:
        _o_sv = 15'b101001101111110;
      12'b111001111011:
        _o_sv = 15'b101001110000011;
      12'b111001111100:
        _o_sv = 15'b101001110001000;
      12'b111001111101:
        _o_sv = 15'b101001110001100;
      12'b111001111110:
        _o_sv = 15'b101001110010001;
      12'b111001111111:
        _o_sv = 15'b101001110010110;
      12'b111010000000:
        _o_sv = 15'b101001110011011;
      12'b111010000001:
        _o_sv = 15'b101001110011111;
      12'b111010000010:
        _o_sv = 15'b101001110100100;
      12'b111010000011:
        _o_sv = 15'b101001110101001;
      12'b111010000100:
        _o_sv = 15'b101001110101110;
      12'b111010000101:
        _o_sv = 15'b101001110110010;
      12'b111010000110:
        _o_sv = 15'b101001110110111;
      12'b111010000111:
        _o_sv = 15'b101001110111100;
      12'b111010001000:
        _o_sv = 15'b101001111000001;
      12'b111010001001:
        _o_sv = 15'b101001111000101;
      12'b111010001010:
        _o_sv = 15'b101001111001010;
      12'b111010001011:
        _o_sv = 15'b101001111001111;
      12'b111010001100:
        _o_sv = 15'b101001111010100;
      12'b111010001101:
        _o_sv = 15'b101001111011000;
      12'b111010001110:
        _o_sv = 15'b101001111011101;
      12'b111010001111:
        _o_sv = 15'b101001111100010;
      12'b111010010000:
        _o_sv = 15'b101001111100111;
      12'b111010010001:
        _o_sv = 15'b101001111101011;
      12'b111010010010:
        _o_sv = 15'b101001111110000;
      12'b111010010011:
        _o_sv = 15'b101001111110101;
      12'b111010010100:
        _o_sv = 15'b101001111111010;
      12'b111010010101:
        _o_sv = 15'b101001111111110;
      12'b111010010110:
        _o_sv = 15'b101010000000011;
      12'b111010010111:
        _o_sv = 15'b101010000001000;
      12'b111010011000:
        _o_sv = 15'b101010000001101;
      12'b111010011001:
        _o_sv = 15'b101010000010001;
      12'b111010011010:
        _o_sv = 15'b101010000010110;
      12'b111010011011:
        _o_sv = 15'b101010000011011;
      12'b111010011100:
        _o_sv = 15'b101010000100000;
      12'b111010011101:
        _o_sv = 15'b101010000100100;
      12'b111010011110:
        _o_sv = 15'b101010000101001;
      12'b111010011111:
        _o_sv = 15'b101010000101110;
      12'b111010100000:
        _o_sv = 15'b101010000110011;
      12'b111010100001:
        _o_sv = 15'b101010000110111;
      12'b111010100010:
        _o_sv = 15'b101010000111100;
      12'b111010100011:
        _o_sv = 15'b101010001000001;
      12'b111010100100:
        _o_sv = 15'b101010001000101;
      12'b111010100101:
        _o_sv = 15'b101010001001010;
      12'b111010100110:
        _o_sv = 15'b101010001001111;
      12'b111010100111:
        _o_sv = 15'b101010001010100;
      12'b111010101000:
        _o_sv = 15'b101010001011000;
      12'b111010101001:
        _o_sv = 15'b101010001011101;
      12'b111010101010:
        _o_sv = 15'b101010001100010;
      12'b111010101011:
        _o_sv = 15'b101010001100111;
      12'b111010101100:
        _o_sv = 15'b101010001101011;
      12'b111010101101:
        _o_sv = 15'b101010001110000;
      12'b111010101110:
        _o_sv = 15'b101010001110101;
      12'b111010101111:
        _o_sv = 15'b101010001111001;
      12'b111010110000:
        _o_sv = 15'b101010001111110;
      12'b111010110001:
        _o_sv = 15'b101010010000011;
      12'b111010110010:
        _o_sv = 15'b101010010001000;
      12'b111010110011:
        _o_sv = 15'b101010010001100;
      12'b111010110100:
        _o_sv = 15'b101010010010001;
      12'b111010110101:
        _o_sv = 15'b101010010010110;
      12'b111010110110:
        _o_sv = 15'b101010010011010;
      12'b111010110111:
        _o_sv = 15'b101010010011111;
      12'b111010111000:
        _o_sv = 15'b101010010100100;
      12'b111010111001:
        _o_sv = 15'b101010010101001;
      12'b111010111010:
        _o_sv = 15'b101010010101101;
      12'b111010111011:
        _o_sv = 15'b101010010110010;
      12'b111010111100:
        _o_sv = 15'b101010010110111;
      12'b111010111101:
        _o_sv = 15'b101010010111011;
      12'b111010111110:
        _o_sv = 15'b101010011000000;
      12'b111010111111:
        _o_sv = 15'b101010011000101;
      12'b111011000000:
        _o_sv = 15'b101010011001010;
      12'b111011000001:
        _o_sv = 15'b101010011001110;
      12'b111011000010:
        _o_sv = 15'b101010011010011;
      12'b111011000011:
        _o_sv = 15'b101010011011000;
      12'b111011000100:
        _o_sv = 15'b101010011011100;
      12'b111011000101:
        _o_sv = 15'b101010011100001;
      12'b111011000110:
        _o_sv = 15'b101010011100110;
      12'b111011000111:
        _o_sv = 15'b101010011101010;
      12'b111011001000:
        _o_sv = 15'b101010011101111;
      12'b111011001001:
        _o_sv = 15'b101010011110100;
      12'b111011001010:
        _o_sv = 15'b101010011111001;
      12'b111011001011:
        _o_sv = 15'b101010011111101;
      12'b111011001100:
        _o_sv = 15'b101010100000010;
      12'b111011001101:
        _o_sv = 15'b101010100000111;
      12'b111011001110:
        _o_sv = 15'b101010100001011;
      12'b111011001111:
        _o_sv = 15'b101010100010000;
      12'b111011010000:
        _o_sv = 15'b101010100010101;
      12'b111011010001:
        _o_sv = 15'b101010100011001;
      12'b111011010010:
        _o_sv = 15'b101010100011110;
      12'b111011010011:
        _o_sv = 15'b101010100100011;
      12'b111011010100:
        _o_sv = 15'b101010100101000;
      12'b111011010101:
        _o_sv = 15'b101010100101100;
      12'b111011010110:
        _o_sv = 15'b101010100110001;
      12'b111011010111:
        _o_sv = 15'b101010100110110;
      12'b111011011000:
        _o_sv = 15'b101010100111010;
      12'b111011011001:
        _o_sv = 15'b101010100111111;
      12'b111011011010:
        _o_sv = 15'b101010101000100;
      12'b111011011011:
        _o_sv = 15'b101010101001000;
      12'b111011011100:
        _o_sv = 15'b101010101001101;
      12'b111011011101:
        _o_sv = 15'b101010101010010;
      12'b111011011110:
        _o_sv = 15'b101010101010110;
      12'b111011011111:
        _o_sv = 15'b101010101011011;
      12'b111011100000:
        _o_sv = 15'b101010101100000;
      12'b111011100001:
        _o_sv = 15'b101010101100100;
      12'b111011100010:
        _o_sv = 15'b101010101101001;
      12'b111011100011:
        _o_sv = 15'b101010101101110;
      12'b111011100100:
        _o_sv = 15'b101010101110010;
      12'b111011100101:
        _o_sv = 15'b101010101110111;
      12'b111011100110:
        _o_sv = 15'b101010101111100;
      12'b111011100111:
        _o_sv = 15'b101010110000001;
      12'b111011101000:
        _o_sv = 15'b101010110000101;
      12'b111011101001:
        _o_sv = 15'b101010110001010;
      12'b111011101010:
        _o_sv = 15'b101010110001111;
      12'b111011101011:
        _o_sv = 15'b101010110010011;
      12'b111011101100:
        _o_sv = 15'b101010110011000;
      12'b111011101101:
        _o_sv = 15'b101010110011101;
      12'b111011101110:
        _o_sv = 15'b101010110100001;
      12'b111011101111:
        _o_sv = 15'b101010110100110;
      12'b111011110000:
        _o_sv = 15'b101010110101011;
      12'b111011110001:
        _o_sv = 15'b101010110101111;
      12'b111011110010:
        _o_sv = 15'b101010110110100;
      12'b111011110011:
        _o_sv = 15'b101010110111001;
      12'b111011110100:
        _o_sv = 15'b101010110111101;
      12'b111011110101:
        _o_sv = 15'b101010111000010;
      12'b111011110110:
        _o_sv = 15'b101010111000111;
      12'b111011110111:
        _o_sv = 15'b101010111001011;
      12'b111011111000:
        _o_sv = 15'b101010111010000;
      12'b111011111001:
        _o_sv = 15'b101010111010101;
      12'b111011111010:
        _o_sv = 15'b101010111011001;
      12'b111011111011:
        _o_sv = 15'b101010111011110;
      12'b111011111100:
        _o_sv = 15'b101010111100011;
      12'b111011111101:
        _o_sv = 15'b101010111100111;
      12'b111011111110:
        _o_sv = 15'b101010111101100;
      12'b111011111111:
        _o_sv = 15'b101010111110000;
      12'b111100000000:
        _o_sv = 15'b101010111110101;
      12'b111100000001:
        _o_sv = 15'b101010111111010;
      12'b111100000010:
        _o_sv = 15'b101010111111110;
      12'b111100000011:
        _o_sv = 15'b101011000000011;
      12'b111100000100:
        _o_sv = 15'b101011000001000;
      12'b111100000101:
        _o_sv = 15'b101011000001100;
      12'b111100000110:
        _o_sv = 15'b101011000010001;
      12'b111100000111:
        _o_sv = 15'b101011000010110;
      12'b111100001000:
        _o_sv = 15'b101011000011010;
      12'b111100001001:
        _o_sv = 15'b101011000011111;
      12'b111100001010:
        _o_sv = 15'b101011000100100;
      12'b111100001011:
        _o_sv = 15'b101011000101000;
      12'b111100001100:
        _o_sv = 15'b101011000101101;
      12'b111100001101:
        _o_sv = 15'b101011000110010;
      12'b111100001110:
        _o_sv = 15'b101011000110110;
      12'b111100001111:
        _o_sv = 15'b101011000111011;
      12'b111100010000:
        _o_sv = 15'b101011001000000;
      12'b111100010001:
        _o_sv = 15'b101011001000100;
      12'b111100010010:
        _o_sv = 15'b101011001001001;
      12'b111100010011:
        _o_sv = 15'b101011001001101;
      12'b111100010100:
        _o_sv = 15'b101011001010010;
      12'b111100010101:
        _o_sv = 15'b101011001010111;
      12'b111100010110:
        _o_sv = 15'b101011001011011;
      12'b111100010111:
        _o_sv = 15'b101011001100000;
      12'b111100011000:
        _o_sv = 15'b101011001100101;
      12'b111100011001:
        _o_sv = 15'b101011001101001;
      12'b111100011010:
        _o_sv = 15'b101011001101110;
      12'b111100011011:
        _o_sv = 15'b101011001110011;
      12'b111100011100:
        _o_sv = 15'b101011001110111;
      12'b111100011101:
        _o_sv = 15'b101011001111100;
      12'b111100011110:
        _o_sv = 15'b101011010000000;
      12'b111100011111:
        _o_sv = 15'b101011010000101;
      12'b111100100000:
        _o_sv = 15'b101011010001010;
      12'b111100100001:
        _o_sv = 15'b101011010001110;
      12'b111100100010:
        _o_sv = 15'b101011010010011;
      12'b111100100011:
        _o_sv = 15'b101011010011000;
      12'b111100100100:
        _o_sv = 15'b101011010011100;
      12'b111100100101:
        _o_sv = 15'b101011010100001;
      12'b111100100110:
        _o_sv = 15'b101011010100101;
      12'b111100100111:
        _o_sv = 15'b101011010101010;
      12'b111100101000:
        _o_sv = 15'b101011010101111;
      12'b111100101001:
        _o_sv = 15'b101011010110011;
      12'b111100101010:
        _o_sv = 15'b101011010111000;
      12'b111100101011:
        _o_sv = 15'b101011010111101;
      12'b111100101100:
        _o_sv = 15'b101011011000001;
      12'b111100101101:
        _o_sv = 15'b101011011000110;
      12'b111100101110:
        _o_sv = 15'b101011011001010;
      12'b111100101111:
        _o_sv = 15'b101011011001111;
      12'b111100110000:
        _o_sv = 15'b101011011010100;
      12'b111100110001:
        _o_sv = 15'b101011011011000;
      12'b111100110010:
        _o_sv = 15'b101011011011101;
      12'b111100110011:
        _o_sv = 15'b101011011100010;
      12'b111100110100:
        _o_sv = 15'b101011011100110;
      12'b111100110101:
        _o_sv = 15'b101011011101011;
      12'b111100110110:
        _o_sv = 15'b101011011101111;
      12'b111100110111:
        _o_sv = 15'b101011011110100;
      12'b111100111000:
        _o_sv = 15'b101011011111001;
      12'b111100111001:
        _o_sv = 15'b101011011111101;
      12'b111100111010:
        _o_sv = 15'b101011100000010;
      12'b111100111011:
        _o_sv = 15'b101011100000110;
      12'b111100111100:
        _o_sv = 15'b101011100001011;
      12'b111100111101:
        _o_sv = 15'b101011100010000;
      12'b111100111110:
        _o_sv = 15'b101011100010100;
      12'b111100111111:
        _o_sv = 15'b101011100011001;
      12'b111101000000:
        _o_sv = 15'b101011100011101;
      12'b111101000001:
        _o_sv = 15'b101011100100010;
      12'b111101000010:
        _o_sv = 15'b101011100100111;
      12'b111101000011:
        _o_sv = 15'b101011100101011;
      12'b111101000100:
        _o_sv = 15'b101011100110000;
      12'b111101000101:
        _o_sv = 15'b101011100110100;
      12'b111101000110:
        _o_sv = 15'b101011100111001;
      12'b111101000111:
        _o_sv = 15'b101011100111110;
      12'b111101001000:
        _o_sv = 15'b101011101000010;
      12'b111101001001:
        _o_sv = 15'b101011101000111;
      12'b111101001010:
        _o_sv = 15'b101011101001011;
      12'b111101001011:
        _o_sv = 15'b101011101010000;
      12'b111101001100:
        _o_sv = 15'b101011101010101;
      12'b111101001101:
        _o_sv = 15'b101011101011001;
      12'b111101001110:
        _o_sv = 15'b101011101011110;
      12'b111101001111:
        _o_sv = 15'b101011101100010;
      12'b111101010000:
        _o_sv = 15'b101011101100111;
      12'b111101010001:
        _o_sv = 15'b101011101101100;
      12'b111101010010:
        _o_sv = 15'b101011101110000;
      12'b111101010011:
        _o_sv = 15'b101011101110101;
      12'b111101010100:
        _o_sv = 15'b101011101111001;
      12'b111101010101:
        _o_sv = 15'b101011101111110;
      12'b111101010110:
        _o_sv = 15'b101011110000011;
      12'b111101010111:
        _o_sv = 15'b101011110000111;
      12'b111101011000:
        _o_sv = 15'b101011110001100;
      12'b111101011001:
        _o_sv = 15'b101011110010000;
      12'b111101011010:
        _o_sv = 15'b101011110010101;
      12'b111101011011:
        _o_sv = 15'b101011110011001;
      12'b111101011100:
        _o_sv = 15'b101011110011110;
      12'b111101011101:
        _o_sv = 15'b101011110100011;
      12'b111101011110:
        _o_sv = 15'b101011110100111;
      12'b111101011111:
        _o_sv = 15'b101011110101100;
      12'b111101100000:
        _o_sv = 15'b101011110110000;
      12'b111101100001:
        _o_sv = 15'b101011110110101;
      12'b111101100010:
        _o_sv = 15'b101011110111001;
      12'b111101100011:
        _o_sv = 15'b101011110111110;
      12'b111101100100:
        _o_sv = 15'b101011111000011;
      12'b111101100101:
        _o_sv = 15'b101011111000111;
      12'b111101100110:
        _o_sv = 15'b101011111001100;
      12'b111101100111:
        _o_sv = 15'b101011111010000;
      12'b111101101000:
        _o_sv = 15'b101011111010101;
      12'b111101101001:
        _o_sv = 15'b101011111011001;
      12'b111101101010:
        _o_sv = 15'b101011111011110;
      12'b111101101011:
        _o_sv = 15'b101011111100011;
      12'b111101101100:
        _o_sv = 15'b101011111100111;
      12'b111101101101:
        _o_sv = 15'b101011111101100;
      12'b111101101110:
        _o_sv = 15'b101011111110000;
      12'b111101101111:
        _o_sv = 15'b101011111110101;
      12'b111101110000:
        _o_sv = 15'b101011111111001;
      12'b111101110001:
        _o_sv = 15'b101011111111110;
      12'b111101110010:
        _o_sv = 15'b101100000000011;
      12'b111101110011:
        _o_sv = 15'b101100000000111;
      12'b111101110100:
        _o_sv = 15'b101100000001100;
      12'b111101110101:
        _o_sv = 15'b101100000010000;
      12'b111101110110:
        _o_sv = 15'b101100000010101;
      12'b111101110111:
        _o_sv = 15'b101100000011001;
      12'b111101111000:
        _o_sv = 15'b101100000011110;
      12'b111101111001:
        _o_sv = 15'b101100000100010;
      12'b111101111010:
        _o_sv = 15'b101100000100111;
      12'b111101111011:
        _o_sv = 15'b101100000101100;
      12'b111101111100:
        _o_sv = 15'b101100000110000;
      12'b111101111101:
        _o_sv = 15'b101100000110101;
      12'b111101111110:
        _o_sv = 15'b101100000111001;
      12'b111101111111:
        _o_sv = 15'b101100000111110;
      12'b111110000000:
        _o_sv = 15'b101100001000010;
      12'b111110000001:
        _o_sv = 15'b101100001000111;
      12'b111110000010:
        _o_sv = 15'b101100001001011;
      12'b111110000011:
        _o_sv = 15'b101100001010000;
      12'b111110000100:
        _o_sv = 15'b101100001010101;
      12'b111110000101:
        _o_sv = 15'b101100001011001;
      12'b111110000110:
        _o_sv = 15'b101100001011110;
      12'b111110000111:
        _o_sv = 15'b101100001100010;
      12'b111110001000:
        _o_sv = 15'b101100001100111;
      12'b111110001001:
        _o_sv = 15'b101100001101011;
      12'b111110001010:
        _o_sv = 15'b101100001110000;
      12'b111110001011:
        _o_sv = 15'b101100001110100;
      12'b111110001100:
        _o_sv = 15'b101100001111001;
      12'b111110001101:
        _o_sv = 15'b101100001111101;
      12'b111110001110:
        _o_sv = 15'b101100010000010;
      12'b111110001111:
        _o_sv = 15'b101100010000111;
      12'b111110010000:
        _o_sv = 15'b101100010001011;
      12'b111110010001:
        _o_sv = 15'b101100010010000;
      12'b111110010010:
        _o_sv = 15'b101100010010100;
      12'b111110010011:
        _o_sv = 15'b101100010011001;
      12'b111110010100:
        _o_sv = 15'b101100010011101;
      12'b111110010101:
        _o_sv = 15'b101100010100010;
      12'b111110010110:
        _o_sv = 15'b101100010100110;
      12'b111110010111:
        _o_sv = 15'b101100010101011;
      12'b111110011000:
        _o_sv = 15'b101100010101111;
      12'b111110011001:
        _o_sv = 15'b101100010110100;
      12'b111110011010:
        _o_sv = 15'b101100010111000;
      12'b111110011011:
        _o_sv = 15'b101100010111101;
      12'b111110011100:
        _o_sv = 15'b101100011000001;
      12'b111110011101:
        _o_sv = 15'b101100011000110;
      12'b111110011110:
        _o_sv = 15'b101100011001011;
      12'b111110011111:
        _o_sv = 15'b101100011001111;
      12'b111110100000:
        _o_sv = 15'b101100011010100;
      12'b111110100001:
        _o_sv = 15'b101100011011000;
      12'b111110100010:
        _o_sv = 15'b101100011011101;
      12'b111110100011:
        _o_sv = 15'b101100011100001;
      12'b111110100100:
        _o_sv = 15'b101100011100110;
      12'b111110100101:
        _o_sv = 15'b101100011101010;
      12'b111110100110:
        _o_sv = 15'b101100011101111;
      12'b111110100111:
        _o_sv = 15'b101100011110011;
      12'b111110101000:
        _o_sv = 15'b101100011111000;
      12'b111110101001:
        _o_sv = 15'b101100011111100;
      12'b111110101010:
        _o_sv = 15'b101100100000001;
      12'b111110101011:
        _o_sv = 15'b101100100000101;
      12'b111110101100:
        _o_sv = 15'b101100100001010;
      12'b111110101101:
        _o_sv = 15'b101100100001110;
      12'b111110101110:
        _o_sv = 15'b101100100010011;
      12'b111110101111:
        _o_sv = 15'b101100100010111;
      12'b111110110000:
        _o_sv = 15'b101100100011100;
      12'b111110110001:
        _o_sv = 15'b101100100100000;
      12'b111110110010:
        _o_sv = 15'b101100100100101;
      12'b111110110011:
        _o_sv = 15'b101100100101001;
      12'b111110110100:
        _o_sv = 15'b101100100101110;
      12'b111110110101:
        _o_sv = 15'b101100100110010;
      12'b111110110110:
        _o_sv = 15'b101100100110111;
      12'b111110110111:
        _o_sv = 15'b101100100111011;
      12'b111110111000:
        _o_sv = 15'b101100101000000;
      12'b111110111001:
        _o_sv = 15'b101100101000100;
      12'b111110111010:
        _o_sv = 15'b101100101001001;
      12'b111110111011:
        _o_sv = 15'b101100101001101;
      12'b111110111100:
        _o_sv = 15'b101100101010010;
      12'b111110111101:
        _o_sv = 15'b101100101010110;
      12'b111110111110:
        _o_sv = 15'b101100101011011;
      12'b111110111111:
        _o_sv = 15'b101100101011111;
      12'b111111000000:
        _o_sv = 15'b101100101100100;
      12'b111111000001:
        _o_sv = 15'b101100101101000;
      12'b111111000010:
        _o_sv = 15'b101100101101101;
      12'b111111000011:
        _o_sv = 15'b101100101110001;
      12'b111111000100:
        _o_sv = 15'b101100101110110;
      12'b111111000101:
        _o_sv = 15'b101100101111010;
      12'b111111000110:
        _o_sv = 15'b101100101111111;
      12'b111111000111:
        _o_sv = 15'b101100110000011;
      12'b111111001000:
        _o_sv = 15'b101100110001000;
      12'b111111001001:
        _o_sv = 15'b101100110001100;
      12'b111111001010:
        _o_sv = 15'b101100110010001;
      12'b111111001011:
        _o_sv = 15'b101100110010101;
      12'b111111001100:
        _o_sv = 15'b101100110011010;
      12'b111111001101:
        _o_sv = 15'b101100110011110;
      12'b111111001110:
        _o_sv = 15'b101100110100011;
      12'b111111001111:
        _o_sv = 15'b101100110100111;
      12'b111111010000:
        _o_sv = 15'b101100110101100;
      12'b111111010001:
        _o_sv = 15'b101100110110000;
      12'b111111010010:
        _o_sv = 15'b101100110110101;
      12'b111111010011:
        _o_sv = 15'b101100110111001;
      12'b111111010100:
        _o_sv = 15'b101100110111110;
      12'b111111010101:
        _o_sv = 15'b101100111000010;
      12'b111111010110:
        _o_sv = 15'b101100111000111;
      12'b111111010111:
        _o_sv = 15'b101100111001011;
      12'b111111011000:
        _o_sv = 15'b101100111010000;
      12'b111111011001:
        _o_sv = 15'b101100111010100;
      12'b111111011010:
        _o_sv = 15'b101100111011001;
      12'b111111011011:
        _o_sv = 15'b101100111011101;
      12'b111111011100:
        _o_sv = 15'b101100111100001;
      12'b111111011101:
        _o_sv = 15'b101100111100110;
      12'b111111011110:
        _o_sv = 15'b101100111101010;
      12'b111111011111:
        _o_sv = 15'b101100111101111;
      12'b111111100000:
        _o_sv = 15'b101100111110011;
      12'b111111100001:
        _o_sv = 15'b101100111111000;
      12'b111111100010:
        _o_sv = 15'b101100111111100;
      12'b111111100011:
        _o_sv = 15'b101101000000001;
      12'b111111100100:
        _o_sv = 15'b101101000000101;
      12'b111111100101:
        _o_sv = 15'b101101000001010;
      12'b111111100110:
        _o_sv = 15'b101101000001110;
      12'b111111100111:
        _o_sv = 15'b101101000010011;
      12'b111111101000:
        _o_sv = 15'b101101000010111;
      12'b111111101001:
        _o_sv = 15'b101101000011100;
      12'b111111101010:
        _o_sv = 15'b101101000100000;
      12'b111111101011:
        _o_sv = 15'b101101000100100;
      12'b111111101100:
        _o_sv = 15'b101101000101001;
      12'b111111101101:
        _o_sv = 15'b101101000101101;
      12'b111111101110:
        _o_sv = 15'b101101000110010;
      12'b111111101111:
        _o_sv = 15'b101101000110110;
      12'b111111110000:
        _o_sv = 15'b101101000111011;
      12'b111111110001:
        _o_sv = 15'b101101000111111;
      12'b111111110010:
        _o_sv = 15'b101101001000100;
      12'b111111110011:
        _o_sv = 15'b101101001001000;
      12'b111111110100:
        _o_sv = 15'b101101001001101;
      12'b111111110101:
        _o_sv = 15'b101101001010001;
      12'b111111110110:
        _o_sv = 15'b101101001010110;
      12'b111111110111:
        _o_sv = 15'b101101001011010;
      12'b111111111000:
        _o_sv = 15'b101101001011110;
      12'b111111111001:
        _o_sv = 15'b101101001100011;
      12'b111111111010:
        _o_sv = 15'b101101001100111;
      12'b111111111011:
        _o_sv = 15'b101101001101100;
      12'b111111111100:
        _o_sv = 15'b101101001110000;
      12'b111111111101:
        _o_sv = 15'b101101001110101;
      12'b111111111110:
        _o_sv = 15'b101101001111001;
      12'b111111111111:
        _o_sv = 15'b101101001111110;
      13'b1000000000000:
        _o_sv = 15'b101101010000010;
      13'b1000000000001:
        _o_sv = 15'b101101010000110;
      13'b1000000000010:
        _o_sv = 15'b101101010001011;
      13'b1000000000011:
        _o_sv = 15'b101101010001111;
      13'b1000000000100:
        _o_sv = 15'b101101010010100;
      13'b1000000000101:
        _o_sv = 15'b101101010011000;
      13'b1000000000110:
        _o_sv = 15'b101101010011101;
      13'b1000000000111:
        _o_sv = 15'b101101010100001;
      13'b1000000001000:
        _o_sv = 15'b101101010100101;
      13'b1000000001001:
        _o_sv = 15'b101101010101010;
      13'b1000000001010:
        _o_sv = 15'b101101010101110;
      13'b1000000001011:
        _o_sv = 15'b101101010110011;
      13'b1000000001100:
        _o_sv = 15'b101101010110111;
      13'b1000000001101:
        _o_sv = 15'b101101010111100;
      13'b1000000001110:
        _o_sv = 15'b101101011000000;
      13'b1000000001111:
        _o_sv = 15'b101101011000101;
      13'b1000000010000:
        _o_sv = 15'b101101011001001;
      13'b1000000010001:
        _o_sv = 15'b101101011001101;
      13'b1000000010010:
        _o_sv = 15'b101101011010010;
      13'b1000000010011:
        _o_sv = 15'b101101011010110;
      13'b1000000010100:
        _o_sv = 15'b101101011011011;
      13'b1000000010101:
        _o_sv = 15'b101101011011111;
      13'b1000000010110:
        _o_sv = 15'b101101011100100;
      13'b1000000010111:
        _o_sv = 15'b101101011101000;
      13'b1000000011000:
        _o_sv = 15'b101101011101100;
      13'b1000000011001:
        _o_sv = 15'b101101011110001;
      13'b1000000011010:
        _o_sv = 15'b101101011110101;
      13'b1000000011011:
        _o_sv = 15'b101101011111010;
      13'b1000000011100:
        _o_sv = 15'b101101011111110;
      13'b1000000011101:
        _o_sv = 15'b101101100000010;
      13'b1000000011110:
        _o_sv = 15'b101101100000111;
      13'b1000000011111:
        _o_sv = 15'b101101100001011;
      13'b1000000100000:
        _o_sv = 15'b101101100010000;
      13'b1000000100001:
        _o_sv = 15'b101101100010100;
      13'b1000000100010:
        _o_sv = 15'b101101100011001;
      13'b1000000100011:
        _o_sv = 15'b101101100011101;
      13'b1000000100100:
        _o_sv = 15'b101101100100001;
      13'b1000000100101:
        _o_sv = 15'b101101100100110;
      13'b1000000100110:
        _o_sv = 15'b101101100101010;
      13'b1000000100111:
        _o_sv = 15'b101101100101111;
      13'b1000000101000:
        _o_sv = 15'b101101100110011;
      13'b1000000101001:
        _o_sv = 15'b101101100110111;
      13'b1000000101010:
        _o_sv = 15'b101101100111100;
      13'b1000000101011:
        _o_sv = 15'b101101101000000;
      13'b1000000101100:
        _o_sv = 15'b101101101000101;
      13'b1000000101101:
        _o_sv = 15'b101101101001001;
      13'b1000000101110:
        _o_sv = 15'b101101101001101;
      13'b1000000101111:
        _o_sv = 15'b101101101010010;
      13'b1000000110000:
        _o_sv = 15'b101101101010110;
      13'b1000000110001:
        _o_sv = 15'b101101101011011;
      13'b1000000110010:
        _o_sv = 15'b101101101011111;
      13'b1000000110011:
        _o_sv = 15'b101101101100011;
      13'b1000000110100:
        _o_sv = 15'b101101101101000;
      13'b1000000110101:
        _o_sv = 15'b101101101101100;
      13'b1000000110110:
        _o_sv = 15'b101101101110001;
      13'b1000000110111:
        _o_sv = 15'b101101101110101;
      13'b1000000111000:
        _o_sv = 15'b101101101111001;
      13'b1000000111001:
        _o_sv = 15'b101101101111110;
      13'b1000000111010:
        _o_sv = 15'b101101110000010;
      13'b1000000111011:
        _o_sv = 15'b101101110000111;
      13'b1000000111100:
        _o_sv = 15'b101101110001011;
      13'b1000000111101:
        _o_sv = 15'b101101110001111;
      13'b1000000111110:
        _o_sv = 15'b101101110010100;
      13'b1000000111111:
        _o_sv = 15'b101101110011000;
      13'b1000001000000:
        _o_sv = 15'b101101110011101;
      13'b1000001000001:
        _o_sv = 15'b101101110100001;
      13'b1000001000010:
        _o_sv = 15'b101101110100101;
      13'b1000001000011:
        _o_sv = 15'b101101110101010;
      13'b1000001000100:
        _o_sv = 15'b101101110101110;
      13'b1000001000101:
        _o_sv = 15'b101101110110010;
      13'b1000001000110:
        _o_sv = 15'b101101110110111;
      13'b1000001000111:
        _o_sv = 15'b101101110111011;
      13'b1000001001000:
        _o_sv = 15'b101101111000000;
      13'b1000001001001:
        _o_sv = 15'b101101111000100;
      13'b1000001001010:
        _o_sv = 15'b101101111001000;
      13'b1000001001011:
        _o_sv = 15'b101101111001101;
      13'b1000001001100:
        _o_sv = 15'b101101111010001;
      13'b1000001001101:
        _o_sv = 15'b101101111010110;
      13'b1000001001110:
        _o_sv = 15'b101101111011010;
      13'b1000001001111:
        _o_sv = 15'b101101111011110;
      13'b1000001010000:
        _o_sv = 15'b101101111100011;
      13'b1000001010001:
        _o_sv = 15'b101101111100111;
      13'b1000001010010:
        _o_sv = 15'b101101111101011;
      13'b1000001010011:
        _o_sv = 15'b101101111110000;
      13'b1000001010100:
        _o_sv = 15'b101101111110100;
      13'b1000001010101:
        _o_sv = 15'b101101111111001;
      13'b1000001010110:
        _o_sv = 15'b101101111111101;
      13'b1000001010111:
        _o_sv = 15'b101110000000001;
      13'b1000001011000:
        _o_sv = 15'b101110000000110;
      13'b1000001011001:
        _o_sv = 15'b101110000001010;
      13'b1000001011010:
        _o_sv = 15'b101110000001110;
      13'b1000001011011:
        _o_sv = 15'b101110000010011;
      13'b1000001011100:
        _o_sv = 15'b101110000010111;
      13'b1000001011101:
        _o_sv = 15'b101110000011011;
      13'b1000001011110:
        _o_sv = 15'b101110000100000;
      13'b1000001011111:
        _o_sv = 15'b101110000100100;
      13'b1000001100000:
        _o_sv = 15'b101110000101001;
      13'b1000001100001:
        _o_sv = 15'b101110000101101;
      13'b1000001100010:
        _o_sv = 15'b101110000110001;
      13'b1000001100011:
        _o_sv = 15'b101110000110110;
      13'b1000001100100:
        _o_sv = 15'b101110000111010;
      13'b1000001100101:
        _o_sv = 15'b101110000111110;
      13'b1000001100110:
        _o_sv = 15'b101110001000011;
      13'b1000001100111:
        _o_sv = 15'b101110001000111;
      13'b1000001101000:
        _o_sv = 15'b101110001001011;
      13'b1000001101001:
        _o_sv = 15'b101110001010000;
      13'b1000001101010:
        _o_sv = 15'b101110001010100;
      13'b1000001101011:
        _o_sv = 15'b101110001011000;
      13'b1000001101100:
        _o_sv = 15'b101110001011101;
      13'b1000001101101:
        _o_sv = 15'b101110001100001;
      13'b1000001101110:
        _o_sv = 15'b101110001100110;
      13'b1000001101111:
        _o_sv = 15'b101110001101010;
      13'b1000001110000:
        _o_sv = 15'b101110001101110;
      13'b1000001110001:
        _o_sv = 15'b101110001110011;
      13'b1000001110010:
        _o_sv = 15'b101110001110111;
      13'b1000001110011:
        _o_sv = 15'b101110001111011;
      13'b1000001110100:
        _o_sv = 15'b101110010000000;
      13'b1000001110101:
        _o_sv = 15'b101110010000100;
      13'b1000001110110:
        _o_sv = 15'b101110010001000;
      13'b1000001110111:
        _o_sv = 15'b101110010001101;
      13'b1000001111000:
        _o_sv = 15'b101110010010001;
      13'b1000001111001:
        _o_sv = 15'b101110010010101;
      13'b1000001111010:
        _o_sv = 15'b101110010011010;
      13'b1000001111011:
        _o_sv = 15'b101110010011110;
      13'b1000001111100:
        _o_sv = 15'b101110010100010;
      13'b1000001111101:
        _o_sv = 15'b101110010100111;
      13'b1000001111110:
        _o_sv = 15'b101110010101011;
      13'b1000001111111:
        _o_sv = 15'b101110010101111;
      13'b1000010000000:
        _o_sv = 15'b101110010110100;
      13'b1000010000001:
        _o_sv = 15'b101110010111000;
      13'b1000010000010:
        _o_sv = 15'b101110010111100;
      13'b1000010000011:
        _o_sv = 15'b101110011000001;
      13'b1000010000100:
        _o_sv = 15'b101110011000101;
      13'b1000010000101:
        _o_sv = 15'b101110011001001;
      13'b1000010000110:
        _o_sv = 15'b101110011001110;
      13'b1000010000111:
        _o_sv = 15'b101110011010010;
      13'b1000010001000:
        _o_sv = 15'b101110011010110;
      13'b1000010001001:
        _o_sv = 15'b101110011011011;
      13'b1000010001010:
        _o_sv = 15'b101110011011111;
      13'b1000010001011:
        _o_sv = 15'b101110011100011;
      13'b1000010001100:
        _o_sv = 15'b101110011101000;
      13'b1000010001101:
        _o_sv = 15'b101110011101100;
      13'b1000010001110:
        _o_sv = 15'b101110011110000;
      13'b1000010001111:
        _o_sv = 15'b101110011110101;
      13'b1000010010000:
        _o_sv = 15'b101110011111001;
      13'b1000010010001:
        _o_sv = 15'b101110011111101;
      13'b1000010010010:
        _o_sv = 15'b101110100000001;
      13'b1000010010011:
        _o_sv = 15'b101110100000110;
      13'b1000010010100:
        _o_sv = 15'b101110100001010;
      13'b1000010010101:
        _o_sv = 15'b101110100001110;
      13'b1000010010110:
        _o_sv = 15'b101110100010011;
      13'b1000010010111:
        _o_sv = 15'b101110100010111;
      13'b1000010011000:
        _o_sv = 15'b101110100011011;
      13'b1000010011001:
        _o_sv = 15'b101110100100000;
      13'b1000010011010:
        _o_sv = 15'b101110100100100;
      13'b1000010011011:
        _o_sv = 15'b101110100101000;
      13'b1000010011100:
        _o_sv = 15'b101110100101101;
      13'b1000010011101:
        _o_sv = 15'b101110100110001;
      13'b1000010011110:
        _o_sv = 15'b101110100110101;
      13'b1000010011111:
        _o_sv = 15'b101110100111010;
      13'b1000010100000:
        _o_sv = 15'b101110100111110;
      13'b1000010100001:
        _o_sv = 15'b101110101000010;
      13'b1000010100010:
        _o_sv = 15'b101110101000110;
      13'b1000010100011:
        _o_sv = 15'b101110101001011;
      13'b1000010100100:
        _o_sv = 15'b101110101001111;
      13'b1000010100101:
        _o_sv = 15'b101110101010011;
      13'b1000010100110:
        _o_sv = 15'b101110101011000;
      13'b1000010100111:
        _o_sv = 15'b101110101011100;
      13'b1000010101000:
        _o_sv = 15'b101110101100000;
      13'b1000010101001:
        _o_sv = 15'b101110101100101;
      13'b1000010101010:
        _o_sv = 15'b101110101101001;
      13'b1000010101011:
        _o_sv = 15'b101110101101101;
      13'b1000010101100:
        _o_sv = 15'b101110101110001;
      13'b1000010101101:
        _o_sv = 15'b101110101110110;
      13'b1000010101110:
        _o_sv = 15'b101110101111010;
      13'b1000010101111:
        _o_sv = 15'b101110101111110;
      13'b1000010110000:
        _o_sv = 15'b101110110000011;
      13'b1000010110001:
        _o_sv = 15'b101110110000111;
      13'b1000010110010:
        _o_sv = 15'b101110110001011;
      13'b1000010110011:
        _o_sv = 15'b101110110001111;
      13'b1000010110100:
        _o_sv = 15'b101110110010100;
      13'b1000010110101:
        _o_sv = 15'b101110110011000;
      13'b1000010110110:
        _o_sv = 15'b101110110011100;
      13'b1000010110111:
        _o_sv = 15'b101110110100001;
      13'b1000010111000:
        _o_sv = 15'b101110110100101;
      13'b1000010111001:
        _o_sv = 15'b101110110101001;
      13'b1000010111010:
        _o_sv = 15'b101110110101101;
      13'b1000010111011:
        _o_sv = 15'b101110110110010;
      13'b1000010111100:
        _o_sv = 15'b101110110110110;
      13'b1000010111101:
        _o_sv = 15'b101110110111010;
      13'b1000010111110:
        _o_sv = 15'b101110110111111;
      13'b1000010111111:
        _o_sv = 15'b101110111000011;
      13'b1000011000000:
        _o_sv = 15'b101110111000111;
      13'b1000011000001:
        _o_sv = 15'b101110111001011;
      13'b1000011000010:
        _o_sv = 15'b101110111010000;
      13'b1000011000011:
        _o_sv = 15'b101110111010100;
      13'b1000011000100:
        _o_sv = 15'b101110111011000;
      13'b1000011000101:
        _o_sv = 15'b101110111011100;
      13'b1000011000110:
        _o_sv = 15'b101110111100001;
      13'b1000011000111:
        _o_sv = 15'b101110111100101;
      13'b1000011001000:
        _o_sv = 15'b101110111101001;
      13'b1000011001001:
        _o_sv = 15'b101110111101110;
      13'b1000011001010:
        _o_sv = 15'b101110111110010;
      13'b1000011001011:
        _o_sv = 15'b101110111110110;
      13'b1000011001100:
        _o_sv = 15'b101110111111010;
      13'b1000011001101:
        _o_sv = 15'b101110111111111;
      13'b1000011001110:
        _o_sv = 15'b101111000000011;
      13'b1000011001111:
        _o_sv = 15'b101111000000111;
      13'b1000011010000:
        _o_sv = 15'b101111000001011;
      13'b1000011010001:
        _o_sv = 15'b101111000010000;
      13'b1000011010010:
        _o_sv = 15'b101111000010100;
      13'b1000011010011:
        _o_sv = 15'b101111000011000;
      13'b1000011010100:
        _o_sv = 15'b101111000011100;
      13'b1000011010101:
        _o_sv = 15'b101111000100001;
      13'b1000011010110:
        _o_sv = 15'b101111000100101;
      13'b1000011010111:
        _o_sv = 15'b101111000101001;
      13'b1000011011000:
        _o_sv = 15'b101111000101101;
      13'b1000011011001:
        _o_sv = 15'b101111000110010;
      13'b1000011011010:
        _o_sv = 15'b101111000110110;
      13'b1000011011011:
        _o_sv = 15'b101111000111010;
      13'b1000011011100:
        _o_sv = 15'b101111000111111;
      13'b1000011011101:
        _o_sv = 15'b101111001000011;
      13'b1000011011110:
        _o_sv = 15'b101111001000111;
      13'b1000011011111:
        _o_sv = 15'b101111001001011;
      13'b1000011100000:
        _o_sv = 15'b101111001010000;
      13'b1000011100001:
        _o_sv = 15'b101111001010100;
      13'b1000011100010:
        _o_sv = 15'b101111001011000;
      13'b1000011100011:
        _o_sv = 15'b101111001011100;
      13'b1000011100100:
        _o_sv = 15'b101111001100000;
      13'b1000011100101:
        _o_sv = 15'b101111001100101;
      13'b1000011100110:
        _o_sv = 15'b101111001101001;
      13'b1000011100111:
        _o_sv = 15'b101111001101101;
      13'b1000011101000:
        _o_sv = 15'b101111001110001;
      13'b1000011101001:
        _o_sv = 15'b101111001110110;
      13'b1000011101010:
        _o_sv = 15'b101111001111010;
      13'b1000011101011:
        _o_sv = 15'b101111001111110;
      13'b1000011101100:
        _o_sv = 15'b101111010000010;
      13'b1000011101101:
        _o_sv = 15'b101111010000111;
      13'b1000011101110:
        _o_sv = 15'b101111010001011;
      13'b1000011101111:
        _o_sv = 15'b101111010001111;
      13'b1000011110000:
        _o_sv = 15'b101111010010011;
      13'b1000011110001:
        _o_sv = 15'b101111010011000;
      13'b1000011110010:
        _o_sv = 15'b101111010011100;
      13'b1000011110011:
        _o_sv = 15'b101111010100000;
      13'b1000011110100:
        _o_sv = 15'b101111010100100;
      13'b1000011110101:
        _o_sv = 15'b101111010101001;
      13'b1000011110110:
        _o_sv = 15'b101111010101101;
      13'b1000011110111:
        _o_sv = 15'b101111010110001;
      13'b1000011111000:
        _o_sv = 15'b101111010110101;
      13'b1000011111001:
        _o_sv = 15'b101111010111001;
      13'b1000011111010:
        _o_sv = 15'b101111010111110;
      13'b1000011111011:
        _o_sv = 15'b101111011000010;
      13'b1000011111100:
        _o_sv = 15'b101111011000110;
      13'b1000011111101:
        _o_sv = 15'b101111011001010;
      13'b1000011111110:
        _o_sv = 15'b101111011001111;
      13'b1000011111111:
        _o_sv = 15'b101111011010011;
      13'b1000100000000:
        _o_sv = 15'b101111011010111;
      13'b1000100000001:
        _o_sv = 15'b101111011011011;
      13'b1000100000010:
        _o_sv = 15'b101111011011111;
      13'b1000100000011:
        _o_sv = 15'b101111011100100;
      13'b1000100000100:
        _o_sv = 15'b101111011101000;
      13'b1000100000101:
        _o_sv = 15'b101111011101100;
      13'b1000100000110:
        _o_sv = 15'b101111011110000;
      13'b1000100000111:
        _o_sv = 15'b101111011110101;
      13'b1000100001000:
        _o_sv = 15'b101111011111001;
      13'b1000100001001:
        _o_sv = 15'b101111011111101;
      13'b1000100001010:
        _o_sv = 15'b101111100000001;
      13'b1000100001011:
        _o_sv = 15'b101111100000101;
      13'b1000100001100:
        _o_sv = 15'b101111100001010;
      13'b1000100001101:
        _o_sv = 15'b101111100001110;
      13'b1000100001110:
        _o_sv = 15'b101111100010010;
      13'b1000100001111:
        _o_sv = 15'b101111100010110;
      13'b1000100010000:
        _o_sv = 15'b101111100011010;
      13'b1000100010001:
        _o_sv = 15'b101111100011111;
      13'b1000100010010:
        _o_sv = 15'b101111100100011;
      13'b1000100010011:
        _o_sv = 15'b101111100100111;
      13'b1000100010100:
        _o_sv = 15'b101111100101011;
      13'b1000100010101:
        _o_sv = 15'b101111100101111;
      13'b1000100010110:
        _o_sv = 15'b101111100110100;
      13'b1000100010111:
        _o_sv = 15'b101111100111000;
      13'b1000100011000:
        _o_sv = 15'b101111100111100;
      13'b1000100011001:
        _o_sv = 15'b101111101000000;
      13'b1000100011010:
        _o_sv = 15'b101111101000100;
      13'b1000100011011:
        _o_sv = 15'b101111101001001;
      13'b1000100011100:
        _o_sv = 15'b101111101001101;
      13'b1000100011101:
        _o_sv = 15'b101111101010001;
      13'b1000100011110:
        _o_sv = 15'b101111101010101;
      13'b1000100011111:
        _o_sv = 15'b101111101011001;
      13'b1000100100000:
        _o_sv = 15'b101111101011110;
      13'b1000100100001:
        _o_sv = 15'b101111101100010;
      13'b1000100100010:
        _o_sv = 15'b101111101100110;
      13'b1000100100011:
        _o_sv = 15'b101111101101010;
      13'b1000100100100:
        _o_sv = 15'b101111101101110;
      13'b1000100100101:
        _o_sv = 15'b101111101110010;
      13'b1000100100110:
        _o_sv = 15'b101111101110111;
      13'b1000100100111:
        _o_sv = 15'b101111101111011;
      13'b1000100101000:
        _o_sv = 15'b101111101111111;
      13'b1000100101001:
        _o_sv = 15'b101111110000011;
      13'b1000100101010:
        _o_sv = 15'b101111110000111;
      13'b1000100101011:
        _o_sv = 15'b101111110001100;
      13'b1000100101100:
        _o_sv = 15'b101111110010000;
      13'b1000100101101:
        _o_sv = 15'b101111110010100;
      13'b1000100101110:
        _o_sv = 15'b101111110011000;
      13'b1000100101111:
        _o_sv = 15'b101111110011100;
      13'b1000100110000:
        _o_sv = 15'b101111110100000;
      13'b1000100110001:
        _o_sv = 15'b101111110100101;
      13'b1000100110010:
        _o_sv = 15'b101111110101001;
      13'b1000100110011:
        _o_sv = 15'b101111110101101;
      13'b1000100110100:
        _o_sv = 15'b101111110110001;
      13'b1000100110101:
        _o_sv = 15'b101111110110101;
      13'b1000100110110:
        _o_sv = 15'b101111110111010;
      13'b1000100110111:
        _o_sv = 15'b101111110111110;
      13'b1000100111000:
        _o_sv = 15'b101111111000010;
      13'b1000100111001:
        _o_sv = 15'b101111111000110;
      13'b1000100111010:
        _o_sv = 15'b101111111001010;
      13'b1000100111011:
        _o_sv = 15'b101111111001110;
      13'b1000100111100:
        _o_sv = 15'b101111111010011;
      13'b1000100111101:
        _o_sv = 15'b101111111010111;
      13'b1000100111110:
        _o_sv = 15'b101111111011011;
      13'b1000100111111:
        _o_sv = 15'b101111111011111;
      13'b1000101000000:
        _o_sv = 15'b101111111100011;
      13'b1000101000001:
        _o_sv = 15'b101111111100111;
      13'b1000101000010:
        _o_sv = 15'b101111111101100;
      13'b1000101000011:
        _o_sv = 15'b101111111110000;
      13'b1000101000100:
        _o_sv = 15'b101111111110100;
      13'b1000101000101:
        _o_sv = 15'b101111111111000;
      13'b1000101000110:
        _o_sv = 15'b101111111111100;
      13'b1000101000111:
        _o_sv = 15'b110000000000000;
      13'b1000101001000:
        _o_sv = 15'b110000000000100;
      13'b1000101001001:
        _o_sv = 15'b110000000001001;
      13'b1000101001010:
        _o_sv = 15'b110000000001101;
      13'b1000101001011:
        _o_sv = 15'b110000000010001;
      13'b1000101001100:
        _o_sv = 15'b110000000010101;
      13'b1000101001101:
        _o_sv = 15'b110000000011001;
      13'b1000101001110:
        _o_sv = 15'b110000000011101;
      13'b1000101001111:
        _o_sv = 15'b110000000100010;
      13'b1000101010000:
        _o_sv = 15'b110000000100110;
      13'b1000101010001:
        _o_sv = 15'b110000000101010;
      13'b1000101010010:
        _o_sv = 15'b110000000101110;
      13'b1000101010011:
        _o_sv = 15'b110000000110010;
      13'b1000101010100:
        _o_sv = 15'b110000000110110;
      13'b1000101010101:
        _o_sv = 15'b110000000111010;
      13'b1000101010110:
        _o_sv = 15'b110000000111111;
      13'b1000101010111:
        _o_sv = 15'b110000001000011;
      13'b1000101011000:
        _o_sv = 15'b110000001000111;
      13'b1000101011001:
        _o_sv = 15'b110000001001011;
      13'b1000101011010:
        _o_sv = 15'b110000001001111;
      13'b1000101011011:
        _o_sv = 15'b110000001010011;
      13'b1000101011100:
        _o_sv = 15'b110000001010111;
      13'b1000101011101:
        _o_sv = 15'b110000001011100;
      13'b1000101011110:
        _o_sv = 15'b110000001100000;
      13'b1000101011111:
        _o_sv = 15'b110000001100100;
      13'b1000101100000:
        _o_sv = 15'b110000001101000;
      13'b1000101100001:
        _o_sv = 15'b110000001101100;
      13'b1000101100010:
        _o_sv = 15'b110000001110000;
      13'b1000101100011:
        _o_sv = 15'b110000001110100;
      13'b1000101100100:
        _o_sv = 15'b110000001111000;
      13'b1000101100101:
        _o_sv = 15'b110000001111101;
      13'b1000101100110:
        _o_sv = 15'b110000010000001;
      13'b1000101100111:
        _o_sv = 15'b110000010000101;
      13'b1000101101000:
        _o_sv = 15'b110000010001001;
      13'b1000101101001:
        _o_sv = 15'b110000010001101;
      13'b1000101101010:
        _o_sv = 15'b110000010010001;
      13'b1000101101011:
        _o_sv = 15'b110000010010101;
      13'b1000101101100:
        _o_sv = 15'b110000010011001;
      13'b1000101101101:
        _o_sv = 15'b110000010011110;
      13'b1000101101110:
        _o_sv = 15'b110000010100010;
      13'b1000101101111:
        _o_sv = 15'b110000010100110;
      13'b1000101110000:
        _o_sv = 15'b110000010101010;
      13'b1000101110001:
        _o_sv = 15'b110000010101110;
      13'b1000101110010:
        _o_sv = 15'b110000010110010;
      13'b1000101110011:
        _o_sv = 15'b110000010110110;
      13'b1000101110100:
        _o_sv = 15'b110000010111010;
      13'b1000101110101:
        _o_sv = 15'b110000010111111;
      13'b1000101110110:
        _o_sv = 15'b110000011000011;
      13'b1000101110111:
        _o_sv = 15'b110000011000111;
      13'b1000101111000:
        _o_sv = 15'b110000011001011;
      13'b1000101111001:
        _o_sv = 15'b110000011001111;
      13'b1000101111010:
        _o_sv = 15'b110000011010011;
      13'b1000101111011:
        _o_sv = 15'b110000011010111;
      13'b1000101111100:
        _o_sv = 15'b110000011011011;
      13'b1000101111101:
        _o_sv = 15'b110000011011111;
      13'b1000101111110:
        _o_sv = 15'b110000011100100;
      13'b1000101111111:
        _o_sv = 15'b110000011101000;
      13'b1000110000000:
        _o_sv = 15'b110000011101100;
      13'b1000110000001:
        _o_sv = 15'b110000011110000;
      13'b1000110000010:
        _o_sv = 15'b110000011110100;
      13'b1000110000011:
        _o_sv = 15'b110000011111000;
      13'b1000110000100:
        _o_sv = 15'b110000011111100;
      13'b1000110000101:
        _o_sv = 15'b110000100000000;
      13'b1000110000110:
        _o_sv = 15'b110000100000100;
      13'b1000110000111:
        _o_sv = 15'b110000100001000;
      13'b1000110001000:
        _o_sv = 15'b110000100001101;
      13'b1000110001001:
        _o_sv = 15'b110000100010001;
      13'b1000110001010:
        _o_sv = 15'b110000100010101;
      13'b1000110001011:
        _o_sv = 15'b110000100011001;
      13'b1000110001100:
        _o_sv = 15'b110000100011101;
      13'b1000110001101:
        _o_sv = 15'b110000100100001;
      13'b1000110001110:
        _o_sv = 15'b110000100100101;
      13'b1000110001111:
        _o_sv = 15'b110000100101001;
      13'b1000110010000:
        _o_sv = 15'b110000100101101;
      13'b1000110010001:
        _o_sv = 15'b110000100110001;
      13'b1000110010010:
        _o_sv = 15'b110000100110101;
      13'b1000110010011:
        _o_sv = 15'b110000100111010;
      13'b1000110010100:
        _o_sv = 15'b110000100111110;
      13'b1000110010101:
        _o_sv = 15'b110000101000010;
      13'b1000110010110:
        _o_sv = 15'b110000101000110;
      13'b1000110010111:
        _o_sv = 15'b110000101001010;
      13'b1000110011000:
        _o_sv = 15'b110000101001110;
      13'b1000110011001:
        _o_sv = 15'b110000101010010;
      13'b1000110011010:
        _o_sv = 15'b110000101010110;
      13'b1000110011011:
        _o_sv = 15'b110000101011010;
      13'b1000110011100:
        _o_sv = 15'b110000101011110;
      13'b1000110011101:
        _o_sv = 15'b110000101100010;
      13'b1000110011110:
        _o_sv = 15'b110000101100110;
      13'b1000110011111:
        _o_sv = 15'b110000101101011;
      13'b1000110100000:
        _o_sv = 15'b110000101101111;
      13'b1000110100001:
        _o_sv = 15'b110000101110011;
      13'b1000110100010:
        _o_sv = 15'b110000101110111;
      13'b1000110100011:
        _o_sv = 15'b110000101111011;
      13'b1000110100100:
        _o_sv = 15'b110000101111111;
      13'b1000110100101:
        _o_sv = 15'b110000110000011;
      13'b1000110100110:
        _o_sv = 15'b110000110000111;
      13'b1000110100111:
        _o_sv = 15'b110000110001011;
      13'b1000110101000:
        _o_sv = 15'b110000110001111;
      13'b1000110101001:
        _o_sv = 15'b110000110010011;
      13'b1000110101010:
        _o_sv = 15'b110000110010111;
      13'b1000110101011:
        _o_sv = 15'b110000110011011;
      13'b1000110101100:
        _o_sv = 15'b110000110011111;
      13'b1000110101101:
        _o_sv = 15'b110000110100011;
      13'b1000110101110:
        _o_sv = 15'b110000110101000;
      13'b1000110101111:
        _o_sv = 15'b110000110101100;
      13'b1000110110000:
        _o_sv = 15'b110000110110000;
      13'b1000110110001:
        _o_sv = 15'b110000110110100;
      13'b1000110110010:
        _o_sv = 15'b110000110111000;
      13'b1000110110011:
        _o_sv = 15'b110000110111100;
      13'b1000110110100:
        _o_sv = 15'b110000111000000;
      13'b1000110110101:
        _o_sv = 15'b110000111000100;
      13'b1000110110110:
        _o_sv = 15'b110000111001000;
      13'b1000110110111:
        _o_sv = 15'b110000111001100;
      13'b1000110111000:
        _o_sv = 15'b110000111010000;
      13'b1000110111001:
        _o_sv = 15'b110000111010100;
      13'b1000110111010:
        _o_sv = 15'b110000111011000;
      13'b1000110111011:
        _o_sv = 15'b110000111011100;
      13'b1000110111100:
        _o_sv = 15'b110000111100000;
      13'b1000110111101:
        _o_sv = 15'b110000111100100;
      13'b1000110111110:
        _o_sv = 15'b110000111101000;
      13'b1000110111111:
        _o_sv = 15'b110000111101100;
      13'b1000111000000:
        _o_sv = 15'b110000111110001;
      13'b1000111000001:
        _o_sv = 15'b110000111110101;
      13'b1000111000010:
        _o_sv = 15'b110000111111001;
      13'b1000111000011:
        _o_sv = 15'b110000111111101;
      13'b1000111000100:
        _o_sv = 15'b110001000000001;
      13'b1000111000101:
        _o_sv = 15'b110001000000101;
      13'b1000111000110:
        _o_sv = 15'b110001000001001;
      13'b1000111000111:
        _o_sv = 15'b110001000001101;
      13'b1000111001000:
        _o_sv = 15'b110001000010001;
      13'b1000111001001:
        _o_sv = 15'b110001000010101;
      13'b1000111001010:
        _o_sv = 15'b110001000011001;
      13'b1000111001011:
        _o_sv = 15'b110001000011101;
      13'b1000111001100:
        _o_sv = 15'b110001000100001;
      13'b1000111001101:
        _o_sv = 15'b110001000100101;
      13'b1000111001110:
        _o_sv = 15'b110001000101001;
      13'b1000111001111:
        _o_sv = 15'b110001000101101;
      13'b1000111010000:
        _o_sv = 15'b110001000110001;
      13'b1000111010001:
        _o_sv = 15'b110001000110101;
      13'b1000111010010:
        _o_sv = 15'b110001000111001;
      13'b1000111010011:
        _o_sv = 15'b110001000111101;
      13'b1000111010100:
        _o_sv = 15'b110001001000001;
      13'b1000111010101:
        _o_sv = 15'b110001001000101;
      13'b1000111010110:
        _o_sv = 15'b110001001001001;
      13'b1000111010111:
        _o_sv = 15'b110001001001101;
      13'b1000111011000:
        _o_sv = 15'b110001001010001;
      13'b1000111011001:
        _o_sv = 15'b110001001010101;
      13'b1000111011010:
        _o_sv = 15'b110001001011001;
      13'b1000111011011:
        _o_sv = 15'b110001001011101;
      13'b1000111011100:
        _o_sv = 15'b110001001100001;
      13'b1000111011101:
        _o_sv = 15'b110001001100101;
      13'b1000111011110:
        _o_sv = 15'b110001001101001;
      13'b1000111011111:
        _o_sv = 15'b110001001101101;
      13'b1000111100000:
        _o_sv = 15'b110001001110001;
      13'b1000111100001:
        _o_sv = 15'b110001001110101;
      13'b1000111100010:
        _o_sv = 15'b110001001111010;
      13'b1000111100011:
        _o_sv = 15'b110001001111110;
      13'b1000111100100:
        _o_sv = 15'b110001010000010;
      13'b1000111100101:
        _o_sv = 15'b110001010000110;
      13'b1000111100110:
        _o_sv = 15'b110001010001010;
      13'b1000111100111:
        _o_sv = 15'b110001010001110;
      13'b1000111101000:
        _o_sv = 15'b110001010010010;
      13'b1000111101001:
        _o_sv = 15'b110001010010110;
      13'b1000111101010:
        _o_sv = 15'b110001010011010;
      13'b1000111101011:
        _o_sv = 15'b110001010011110;
      13'b1000111101100:
        _o_sv = 15'b110001010100010;
      13'b1000111101101:
        _o_sv = 15'b110001010100110;
      13'b1000111101110:
        _o_sv = 15'b110001010101010;
      13'b1000111101111:
        _o_sv = 15'b110001010101110;
      13'b1000111110000:
        _o_sv = 15'b110001010110010;
      13'b1000111110001:
        _o_sv = 15'b110001010110110;
      13'b1000111110010:
        _o_sv = 15'b110001010111010;
      13'b1000111110011:
        _o_sv = 15'b110001010111110;
      13'b1000111110100:
        _o_sv = 15'b110001011000010;
      13'b1000111110101:
        _o_sv = 15'b110001011000110;
      13'b1000111110110:
        _o_sv = 15'b110001011001010;
      13'b1000111110111:
        _o_sv = 15'b110001011001110;
      13'b1000111111000:
        _o_sv = 15'b110001011010010;
      13'b1000111111001:
        _o_sv = 15'b110001011010110;
      13'b1000111111010:
        _o_sv = 15'b110001011011010;
      13'b1000111111011:
        _o_sv = 15'b110001011011110;
      13'b1000111111100:
        _o_sv = 15'b110001011100010;
      13'b1000111111101:
        _o_sv = 15'b110001011100110;
      13'b1000111111110:
        _o_sv = 15'b110001011101010;
      13'b1000111111111:
        _o_sv = 15'b110001011101110;
      13'b1001000000000:
        _o_sv = 15'b110001011110010;
      13'b1001000000001:
        _o_sv = 15'b110001011110101;
      13'b1001000000010:
        _o_sv = 15'b110001011111001;
      13'b1001000000011:
        _o_sv = 15'b110001011111101;
      13'b1001000000100:
        _o_sv = 15'b110001100000001;
      13'b1001000000101:
        _o_sv = 15'b110001100000101;
      13'b1001000000110:
        _o_sv = 15'b110001100001001;
      13'b1001000000111:
        _o_sv = 15'b110001100001101;
      13'b1001000001000:
        _o_sv = 15'b110001100010001;
      13'b1001000001001:
        _o_sv = 15'b110001100010101;
      13'b1001000001010:
        _o_sv = 15'b110001100011001;
      13'b1001000001011:
        _o_sv = 15'b110001100011101;
      13'b1001000001100:
        _o_sv = 15'b110001100100001;
      13'b1001000001101:
        _o_sv = 15'b110001100100101;
      13'b1001000001110:
        _o_sv = 15'b110001100101001;
      13'b1001000001111:
        _o_sv = 15'b110001100101101;
      13'b1001000010000:
        _o_sv = 15'b110001100110001;
      13'b1001000010001:
        _o_sv = 15'b110001100110101;
      13'b1001000010010:
        _o_sv = 15'b110001100111001;
      13'b1001000010011:
        _o_sv = 15'b110001100111101;
      13'b1001000010100:
        _o_sv = 15'b110001101000001;
      13'b1001000010101:
        _o_sv = 15'b110001101000101;
      13'b1001000010110:
        _o_sv = 15'b110001101001001;
      13'b1001000010111:
        _o_sv = 15'b110001101001101;
      13'b1001000011000:
        _o_sv = 15'b110001101010001;
      13'b1001000011001:
        _o_sv = 15'b110001101010101;
      13'b1001000011010:
        _o_sv = 15'b110001101011001;
      13'b1001000011011:
        _o_sv = 15'b110001101011101;
      13'b1001000011100:
        _o_sv = 15'b110001101100001;
      13'b1001000011101:
        _o_sv = 15'b110001101100101;
      13'b1001000011110:
        _o_sv = 15'b110001101101001;
      13'b1001000011111:
        _o_sv = 15'b110001101101101;
      13'b1001000100000:
        _o_sv = 15'b110001101110001;
      13'b1001000100001:
        _o_sv = 15'b110001101110101;
      13'b1001000100010:
        _o_sv = 15'b110001101111000;
      13'b1001000100011:
        _o_sv = 15'b110001101111100;
      13'b1001000100100:
        _o_sv = 15'b110001110000000;
      13'b1001000100101:
        _o_sv = 15'b110001110000100;
      13'b1001000100110:
        _o_sv = 15'b110001110001000;
      13'b1001000100111:
        _o_sv = 15'b110001110001100;
      13'b1001000101000:
        _o_sv = 15'b110001110010000;
      13'b1001000101001:
        _o_sv = 15'b110001110010100;
      13'b1001000101010:
        _o_sv = 15'b110001110011000;
      13'b1001000101011:
        _o_sv = 15'b110001110011100;
      13'b1001000101100:
        _o_sv = 15'b110001110100000;
      13'b1001000101101:
        _o_sv = 15'b110001110100100;
      13'b1001000101110:
        _o_sv = 15'b110001110101000;
      13'b1001000101111:
        _o_sv = 15'b110001110101100;
      13'b1001000110000:
        _o_sv = 15'b110001110110000;
      13'b1001000110001:
        _o_sv = 15'b110001110110100;
      13'b1001000110010:
        _o_sv = 15'b110001110111000;
      13'b1001000110011:
        _o_sv = 15'b110001110111100;
      13'b1001000110100:
        _o_sv = 15'b110001111000000;
      13'b1001000110101:
        _o_sv = 15'b110001111000011;
      13'b1001000110110:
        _o_sv = 15'b110001111000111;
      13'b1001000110111:
        _o_sv = 15'b110001111001011;
      13'b1001000111000:
        _o_sv = 15'b110001111001111;
      13'b1001000111001:
        _o_sv = 15'b110001111010011;
      13'b1001000111010:
        _o_sv = 15'b110001111010111;
      13'b1001000111011:
        _o_sv = 15'b110001111011011;
      13'b1001000111100:
        _o_sv = 15'b110001111011111;
      13'b1001000111101:
        _o_sv = 15'b110001111100011;
      13'b1001000111110:
        _o_sv = 15'b110001111100111;
      13'b1001000111111:
        _o_sv = 15'b110001111101011;
      13'b1001001000000:
        _o_sv = 15'b110001111101111;
      13'b1001001000001:
        _o_sv = 15'b110001111110011;
      13'b1001001000010:
        _o_sv = 15'b110001111110111;
      13'b1001001000011:
        _o_sv = 15'b110001111111010;
      13'b1001001000100:
        _o_sv = 15'b110001111111110;
      13'b1001001000101:
        _o_sv = 15'b110010000000010;
      13'b1001001000110:
        _o_sv = 15'b110010000000110;
      13'b1001001000111:
        _o_sv = 15'b110010000001010;
      13'b1001001001000:
        _o_sv = 15'b110010000001110;
      13'b1001001001001:
        _o_sv = 15'b110010000010010;
      13'b1001001001010:
        _o_sv = 15'b110010000010110;
      13'b1001001001011:
        _o_sv = 15'b110010000011010;
      13'b1001001001100:
        _o_sv = 15'b110010000011110;
      13'b1001001001101:
        _o_sv = 15'b110010000100010;
      13'b1001001001110:
        _o_sv = 15'b110010000100110;
      13'b1001001001111:
        _o_sv = 15'b110010000101001;
      13'b1001001010000:
        _o_sv = 15'b110010000101101;
      13'b1001001010001:
        _o_sv = 15'b110010000110001;
      13'b1001001010010:
        _o_sv = 15'b110010000110101;
      13'b1001001010011:
        _o_sv = 15'b110010000111001;
      13'b1001001010100:
        _o_sv = 15'b110010000111101;
      13'b1001001010101:
        _o_sv = 15'b110010001000001;
      13'b1001001010110:
        _o_sv = 15'b110010001000101;
      13'b1001001010111:
        _o_sv = 15'b110010001001001;
      13'b1001001011000:
        _o_sv = 15'b110010001001101;
      13'b1001001011001:
        _o_sv = 15'b110010001010001;
      13'b1001001011010:
        _o_sv = 15'b110010001010100;
      13'b1001001011011:
        _o_sv = 15'b110010001011000;
      13'b1001001011100:
        _o_sv = 15'b110010001011100;
      13'b1001001011101:
        _o_sv = 15'b110010001100000;
      13'b1001001011110:
        _o_sv = 15'b110010001100100;
      13'b1001001011111:
        _o_sv = 15'b110010001101000;
      13'b1001001100000:
        _o_sv = 15'b110010001101100;
      13'b1001001100001:
        _o_sv = 15'b110010001110000;
      13'b1001001100010:
        _o_sv = 15'b110010001110100;
      13'b1001001100011:
        _o_sv = 15'b110010001111000;
      13'b1001001100100:
        _o_sv = 15'b110010001111011;
      13'b1001001100101:
        _o_sv = 15'b110010001111111;
      13'b1001001100110:
        _o_sv = 15'b110010010000011;
      13'b1001001100111:
        _o_sv = 15'b110010010000111;
      13'b1001001101000:
        _o_sv = 15'b110010010001011;
      13'b1001001101001:
        _o_sv = 15'b110010010001111;
      13'b1001001101010:
        _o_sv = 15'b110010010010011;
      13'b1001001101011:
        _o_sv = 15'b110010010010111;
      13'b1001001101100:
        _o_sv = 15'b110010010011011;
      13'b1001001101101:
        _o_sv = 15'b110010010011110;
      13'b1001001101110:
        _o_sv = 15'b110010010100010;
      13'b1001001101111:
        _o_sv = 15'b110010010100110;
      13'b1001001110000:
        _o_sv = 15'b110010010101010;
      13'b1001001110001:
        _o_sv = 15'b110010010101110;
      13'b1001001110010:
        _o_sv = 15'b110010010110010;
      13'b1001001110011:
        _o_sv = 15'b110010010110110;
      13'b1001001110100:
        _o_sv = 15'b110010010111010;
      13'b1001001110101:
        _o_sv = 15'b110010010111101;
      13'b1001001110110:
        _o_sv = 15'b110010011000001;
      13'b1001001110111:
        _o_sv = 15'b110010011000101;
      13'b1001001111000:
        _o_sv = 15'b110010011001001;
      13'b1001001111001:
        _o_sv = 15'b110010011001101;
      13'b1001001111010:
        _o_sv = 15'b110010011010001;
      13'b1001001111011:
        _o_sv = 15'b110010011010101;
      13'b1001001111100:
        _o_sv = 15'b110010011011001;
      13'b1001001111101:
        _o_sv = 15'b110010011011100;
      13'b1001001111110:
        _o_sv = 15'b110010011100000;
      13'b1001001111111:
        _o_sv = 15'b110010011100100;
      13'b1001010000000:
        _o_sv = 15'b110010011101000;
      13'b1001010000001:
        _o_sv = 15'b110010011101100;
      13'b1001010000010:
        _o_sv = 15'b110010011110000;
      13'b1001010000011:
        _o_sv = 15'b110010011110100;
      13'b1001010000100:
        _o_sv = 15'b110010011110111;
      13'b1001010000101:
        _o_sv = 15'b110010011111011;
      13'b1001010000110:
        _o_sv = 15'b110010011111111;
      13'b1001010000111:
        _o_sv = 15'b110010100000011;
      13'b1001010001000:
        _o_sv = 15'b110010100000111;
      13'b1001010001001:
        _o_sv = 15'b110010100001011;
      13'b1001010001010:
        _o_sv = 15'b110010100001111;
      13'b1001010001011:
        _o_sv = 15'b110010100010011;
      13'b1001010001100:
        _o_sv = 15'b110010100010110;
      13'b1001010001101:
        _o_sv = 15'b110010100011010;
      13'b1001010001110:
        _o_sv = 15'b110010100011110;
      13'b1001010001111:
        _o_sv = 15'b110010100100010;
      13'b1001010010000:
        _o_sv = 15'b110010100100110;
      13'b1001010010001:
        _o_sv = 15'b110010100101010;
      13'b1001010010010:
        _o_sv = 15'b110010100101101;
      13'b1001010010011:
        _o_sv = 15'b110010100110001;
      13'b1001010010100:
        _o_sv = 15'b110010100110101;
      13'b1001010010101:
        _o_sv = 15'b110010100111001;
      13'b1001010010110:
        _o_sv = 15'b110010100111101;
      13'b1001010010111:
        _o_sv = 15'b110010101000001;
      13'b1001010011000:
        _o_sv = 15'b110010101000101;
      13'b1001010011001:
        _o_sv = 15'b110010101001000;
      13'b1001010011010:
        _o_sv = 15'b110010101001100;
      13'b1001010011011:
        _o_sv = 15'b110010101010000;
      13'b1001010011100:
        _o_sv = 15'b110010101010100;
      13'b1001010011101:
        _o_sv = 15'b110010101011000;
      13'b1001010011110:
        _o_sv = 15'b110010101011100;
      13'b1001010011111:
        _o_sv = 15'b110010101011111;
      13'b1001010100000:
        _o_sv = 15'b110010101100011;
      13'b1001010100001:
        _o_sv = 15'b110010101100111;
      13'b1001010100010:
        _o_sv = 15'b110010101101011;
      13'b1001010100011:
        _o_sv = 15'b110010101101111;
      13'b1001010100100:
        _o_sv = 15'b110010101110011;
      13'b1001010100101:
        _o_sv = 15'b110010101110110;
      13'b1001010100110:
        _o_sv = 15'b110010101111010;
      13'b1001010100111:
        _o_sv = 15'b110010101111110;
      13'b1001010101000:
        _o_sv = 15'b110010110000010;
      13'b1001010101001:
        _o_sv = 15'b110010110000110;
      13'b1001010101010:
        _o_sv = 15'b110010110001010;
      13'b1001010101011:
        _o_sv = 15'b110010110001101;
      13'b1001010101100:
        _o_sv = 15'b110010110010001;
      13'b1001010101101:
        _o_sv = 15'b110010110010101;
      13'b1001010101110:
        _o_sv = 15'b110010110011001;
      13'b1001010101111:
        _o_sv = 15'b110010110011101;
      13'b1001010110000:
        _o_sv = 15'b110010110100000;
      13'b1001010110001:
        _o_sv = 15'b110010110100100;
      13'b1001010110010:
        _o_sv = 15'b110010110101000;
      13'b1001010110011:
        _o_sv = 15'b110010110101100;
      13'b1001010110100:
        _o_sv = 15'b110010110110000;
      13'b1001010110101:
        _o_sv = 15'b110010110110100;
      13'b1001010110110:
        _o_sv = 15'b110010110110111;
      13'b1001010110111:
        _o_sv = 15'b110010110111011;
      13'b1001010111000:
        _o_sv = 15'b110010110111111;
      13'b1001010111001:
        _o_sv = 15'b110010111000011;
      13'b1001010111010:
        _o_sv = 15'b110010111000111;
      13'b1001010111011:
        _o_sv = 15'b110010111001010;
      13'b1001010111100:
        _o_sv = 15'b110010111001110;
      13'b1001010111101:
        _o_sv = 15'b110010111010010;
      13'b1001010111110:
        _o_sv = 15'b110010111010110;
      13'b1001010111111:
        _o_sv = 15'b110010111011010;
      13'b1001011000000:
        _o_sv = 15'b110010111011101;
      13'b1001011000001:
        _o_sv = 15'b110010111100001;
      13'b1001011000010:
        _o_sv = 15'b110010111100101;
      13'b1001011000011:
        _o_sv = 15'b110010111101001;
      13'b1001011000100:
        _o_sv = 15'b110010111101101;
      13'b1001011000101:
        _o_sv = 15'b110010111110000;
      13'b1001011000110:
        _o_sv = 15'b110010111110100;
      13'b1001011000111:
        _o_sv = 15'b110010111111000;
      13'b1001011001000:
        _o_sv = 15'b110010111111100;
      13'b1001011001001:
        _o_sv = 15'b110011000000000;
      13'b1001011001010:
        _o_sv = 15'b110011000000011;
      13'b1001011001011:
        _o_sv = 15'b110011000000111;
      13'b1001011001100:
        _o_sv = 15'b110011000001011;
      13'b1001011001101:
        _o_sv = 15'b110011000001111;
      13'b1001011001110:
        _o_sv = 15'b110011000010011;
      13'b1001011001111:
        _o_sv = 15'b110011000010110;
      13'b1001011010000:
        _o_sv = 15'b110011000011010;
      13'b1001011010001:
        _o_sv = 15'b110011000011110;
      13'b1001011010010:
        _o_sv = 15'b110011000100010;
      13'b1001011010011:
        _o_sv = 15'b110011000100110;
      13'b1001011010100:
        _o_sv = 15'b110011000101001;
      13'b1001011010101:
        _o_sv = 15'b110011000101101;
      13'b1001011010110:
        _o_sv = 15'b110011000110001;
      13'b1001011010111:
        _o_sv = 15'b110011000110101;
      13'b1001011011000:
        _o_sv = 15'b110011000111001;
      13'b1001011011001:
        _o_sv = 15'b110011000111100;
      13'b1001011011010:
        _o_sv = 15'b110011001000000;
      13'b1001011011011:
        _o_sv = 15'b110011001000100;
      13'b1001011011100:
        _o_sv = 15'b110011001001000;
      13'b1001011011101:
        _o_sv = 15'b110011001001011;
      13'b1001011011110:
        _o_sv = 15'b110011001001111;
      13'b1001011011111:
        _o_sv = 15'b110011001010011;
      13'b1001011100000:
        _o_sv = 15'b110011001010111;
      13'b1001011100001:
        _o_sv = 15'b110011001011011;
      13'b1001011100010:
        _o_sv = 15'b110011001011110;
      13'b1001011100011:
        _o_sv = 15'b110011001100010;
      13'b1001011100100:
        _o_sv = 15'b110011001100110;
      13'b1001011100101:
        _o_sv = 15'b110011001101010;
      13'b1001011100110:
        _o_sv = 15'b110011001101101;
      13'b1001011100111:
        _o_sv = 15'b110011001110001;
      13'b1001011101000:
        _o_sv = 15'b110011001110101;
      13'b1001011101001:
        _o_sv = 15'b110011001111001;
      13'b1001011101010:
        _o_sv = 15'b110011001111100;
      13'b1001011101011:
        _o_sv = 15'b110011010000000;
      13'b1001011101100:
        _o_sv = 15'b110011010000100;
      13'b1001011101101:
        _o_sv = 15'b110011010001000;
      13'b1001011101110:
        _o_sv = 15'b110011010001011;
      13'b1001011101111:
        _o_sv = 15'b110011010001111;
      13'b1001011110000:
        _o_sv = 15'b110011010010011;
      13'b1001011110001:
        _o_sv = 15'b110011010010111;
      13'b1001011110010:
        _o_sv = 15'b110011010011011;
      13'b1001011110011:
        _o_sv = 15'b110011010011110;
      13'b1001011110100:
        _o_sv = 15'b110011010100010;
      13'b1001011110101:
        _o_sv = 15'b110011010100110;
      13'b1001011110110:
        _o_sv = 15'b110011010101010;
      13'b1001011110111:
        _o_sv = 15'b110011010101101;
      13'b1001011111000:
        _o_sv = 15'b110011010110001;
      13'b1001011111001:
        _o_sv = 15'b110011010110101;
      13'b1001011111010:
        _o_sv = 15'b110011010111001;
      13'b1001011111011:
        _o_sv = 15'b110011010111100;
      13'b1001011111100:
        _o_sv = 15'b110011011000000;
      13'b1001011111101:
        _o_sv = 15'b110011011000100;
      13'b1001011111110:
        _o_sv = 15'b110011011001000;
      13'b1001011111111:
        _o_sv = 15'b110011011001011;
      13'b1001100000000:
        _o_sv = 15'b110011011001111;
      13'b1001100000001:
        _o_sv = 15'b110011011010011;
      13'b1001100000010:
        _o_sv = 15'b110011011010110;
      13'b1001100000011:
        _o_sv = 15'b110011011011010;
      13'b1001100000100:
        _o_sv = 15'b110011011011110;
      13'b1001100000101:
        _o_sv = 15'b110011011100010;
      13'b1001100000110:
        _o_sv = 15'b110011011100101;
      13'b1001100000111:
        _o_sv = 15'b110011011101001;
      13'b1001100001000:
        _o_sv = 15'b110011011101101;
      13'b1001100001001:
        _o_sv = 15'b110011011110001;
      13'b1001100001010:
        _o_sv = 15'b110011011110100;
      13'b1001100001011:
        _o_sv = 15'b110011011111000;
      13'b1001100001100:
        _o_sv = 15'b110011011111100;
      13'b1001100001101:
        _o_sv = 15'b110011100000000;
      13'b1001100001110:
        _o_sv = 15'b110011100000011;
      13'b1001100001111:
        _o_sv = 15'b110011100000111;
      13'b1001100010000:
        _o_sv = 15'b110011100001011;
      13'b1001100010001:
        _o_sv = 15'b110011100001110;
      13'b1001100010010:
        _o_sv = 15'b110011100010010;
      13'b1001100010011:
        _o_sv = 15'b110011100010110;
      13'b1001100010100:
        _o_sv = 15'b110011100011010;
      13'b1001100010101:
        _o_sv = 15'b110011100011101;
      13'b1001100010110:
        _o_sv = 15'b110011100100001;
      13'b1001100010111:
        _o_sv = 15'b110011100100101;
      13'b1001100011000:
        _o_sv = 15'b110011100101001;
      13'b1001100011001:
        _o_sv = 15'b110011100101100;
      13'b1001100011010:
        _o_sv = 15'b110011100110000;
      13'b1001100011011:
        _o_sv = 15'b110011100110100;
      13'b1001100011100:
        _o_sv = 15'b110011100110111;
      13'b1001100011101:
        _o_sv = 15'b110011100111011;
      13'b1001100011110:
        _o_sv = 15'b110011100111111;
      13'b1001100011111:
        _o_sv = 15'b110011101000011;
      13'b1001100100000:
        _o_sv = 15'b110011101000110;
      13'b1001100100001:
        _o_sv = 15'b110011101001010;
      13'b1001100100010:
        _o_sv = 15'b110011101001110;
      13'b1001100100011:
        _o_sv = 15'b110011101010001;
      13'b1001100100100:
        _o_sv = 15'b110011101010101;
      13'b1001100100101:
        _o_sv = 15'b110011101011001;
      13'b1001100100110:
        _o_sv = 15'b110011101011101;
      13'b1001100100111:
        _o_sv = 15'b110011101100000;
      13'b1001100101000:
        _o_sv = 15'b110011101100100;
      13'b1001100101001:
        _o_sv = 15'b110011101101000;
      13'b1001100101010:
        _o_sv = 15'b110011101101011;
      13'b1001100101011:
        _o_sv = 15'b110011101101111;
      13'b1001100101100:
        _o_sv = 15'b110011101110011;
      13'b1001100101101:
        _o_sv = 15'b110011101110110;
      13'b1001100101110:
        _o_sv = 15'b110011101111010;
      13'b1001100101111:
        _o_sv = 15'b110011101111110;
      13'b1001100110000:
        _o_sv = 15'b110011110000010;
      13'b1001100110001:
        _o_sv = 15'b110011110000101;
      13'b1001100110010:
        _o_sv = 15'b110011110001001;
      13'b1001100110011:
        _o_sv = 15'b110011110001101;
      13'b1001100110100:
        _o_sv = 15'b110011110010000;
      13'b1001100110101:
        _o_sv = 15'b110011110010100;
      13'b1001100110110:
        _o_sv = 15'b110011110011000;
      13'b1001100110111:
        _o_sv = 15'b110011110011011;
      13'b1001100111000:
        _o_sv = 15'b110011110011111;
      13'b1001100111001:
        _o_sv = 15'b110011110100011;
      13'b1001100111010:
        _o_sv = 15'b110011110100110;
      13'b1001100111011:
        _o_sv = 15'b110011110101010;
      13'b1001100111100:
        _o_sv = 15'b110011110101110;
      13'b1001100111101:
        _o_sv = 15'b110011110110010;
      13'b1001100111110:
        _o_sv = 15'b110011110110101;
      13'b1001100111111:
        _o_sv = 15'b110011110111001;
      13'b1001101000000:
        _o_sv = 15'b110011110111101;
      13'b1001101000001:
        _o_sv = 15'b110011111000000;
      13'b1001101000010:
        _o_sv = 15'b110011111000100;
      13'b1001101000011:
        _o_sv = 15'b110011111001000;
      13'b1001101000100:
        _o_sv = 15'b110011111001011;
      13'b1001101000101:
        _o_sv = 15'b110011111001111;
      13'b1001101000110:
        _o_sv = 15'b110011111010011;
      13'b1001101000111:
        _o_sv = 15'b110011111010110;
      13'b1001101001000:
        _o_sv = 15'b110011111011010;
      13'b1001101001001:
        _o_sv = 15'b110011111011110;
      13'b1001101001010:
        _o_sv = 15'b110011111100001;
      13'b1001101001011:
        _o_sv = 15'b110011111100101;
      13'b1001101001100:
        _o_sv = 15'b110011111101001;
      13'b1001101001101:
        _o_sv = 15'b110011111101100;
      13'b1001101001110:
        _o_sv = 15'b110011111110000;
      13'b1001101001111:
        _o_sv = 15'b110011111110100;
      13'b1001101010000:
        _o_sv = 15'b110011111110111;
      13'b1001101010001:
        _o_sv = 15'b110011111111011;
      13'b1001101010010:
        _o_sv = 15'b110011111111111;
      13'b1001101010011:
        _o_sv = 15'b110100000000010;
      13'b1001101010100:
        _o_sv = 15'b110100000000110;
      13'b1001101010101:
        _o_sv = 15'b110100000001010;
      13'b1001101010110:
        _o_sv = 15'b110100000001101;
      13'b1001101010111:
        _o_sv = 15'b110100000010001;
      13'b1001101011000:
        _o_sv = 15'b110100000010101;
      13'b1001101011001:
        _o_sv = 15'b110100000011000;
      13'b1001101011010:
        _o_sv = 15'b110100000011100;
      13'b1001101011011:
        _o_sv = 15'b110100000100000;
      13'b1001101011100:
        _o_sv = 15'b110100000100011;
      13'b1001101011101:
        _o_sv = 15'b110100000100111;
      13'b1001101011110:
        _o_sv = 15'b110100000101011;
      13'b1001101011111:
        _o_sv = 15'b110100000101110;
      13'b1001101100000:
        _o_sv = 15'b110100000110010;
      13'b1001101100001:
        _o_sv = 15'b110100000110101;
      13'b1001101100010:
        _o_sv = 15'b110100000111001;
      13'b1001101100011:
        _o_sv = 15'b110100000111101;
      13'b1001101100100:
        _o_sv = 15'b110100001000000;
      13'b1001101100101:
        _o_sv = 15'b110100001000100;
      13'b1001101100110:
        _o_sv = 15'b110100001001000;
      13'b1001101100111:
        _o_sv = 15'b110100001001011;
      13'b1001101101000:
        _o_sv = 15'b110100001001111;
      13'b1001101101001:
        _o_sv = 15'b110100001010011;
      13'b1001101101010:
        _o_sv = 15'b110100001010110;
      13'b1001101101011:
        _o_sv = 15'b110100001011010;
      13'b1001101101100:
        _o_sv = 15'b110100001011110;
      13'b1001101101101:
        _o_sv = 15'b110100001100001;
      13'b1001101101110:
        _o_sv = 15'b110100001100101;
      13'b1001101101111:
        _o_sv = 15'b110100001101000;
      13'b1001101110000:
        _o_sv = 15'b110100001101100;
      13'b1001101110001:
        _o_sv = 15'b110100001110000;
      13'b1001101110010:
        _o_sv = 15'b110100001110011;
      13'b1001101110011:
        _o_sv = 15'b110100001110111;
      13'b1001101110100:
        _o_sv = 15'b110100001111011;
      13'b1001101110101:
        _o_sv = 15'b110100001111110;
      13'b1001101110110:
        _o_sv = 15'b110100010000010;
      13'b1001101110111:
        _o_sv = 15'b110100010000110;
      13'b1001101111000:
        _o_sv = 15'b110100010001001;
      13'b1001101111001:
        _o_sv = 15'b110100010001101;
      13'b1001101111010:
        _o_sv = 15'b110100010010000;
      13'b1001101111011:
        _o_sv = 15'b110100010010100;
      13'b1001101111100:
        _o_sv = 15'b110100010011000;
      13'b1001101111101:
        _o_sv = 15'b110100010011011;
      13'b1001101111110:
        _o_sv = 15'b110100010011111;
      13'b1001101111111:
        _o_sv = 15'b110100010100011;
      13'b1001110000000:
        _o_sv = 15'b110100010100110;
      13'b1001110000001:
        _o_sv = 15'b110100010101010;
      13'b1001110000010:
        _o_sv = 15'b110100010101101;
      13'b1001110000011:
        _o_sv = 15'b110100010110001;
      13'b1001110000100:
        _o_sv = 15'b110100010110101;
      13'b1001110000101:
        _o_sv = 15'b110100010111000;
      13'b1001110000110:
        _o_sv = 15'b110100010111100;
      13'b1001110000111:
        _o_sv = 15'b110100010111111;
      13'b1001110001000:
        _o_sv = 15'b110100011000011;
      13'b1001110001001:
        _o_sv = 15'b110100011000111;
      13'b1001110001010:
        _o_sv = 15'b110100011001010;
      13'b1001110001011:
        _o_sv = 15'b110100011001110;
      13'b1001110001100:
        _o_sv = 15'b110100011010001;
      13'b1001110001101:
        _o_sv = 15'b110100011010101;
      13'b1001110001110:
        _o_sv = 15'b110100011011001;
      13'b1001110001111:
        _o_sv = 15'b110100011011100;
      13'b1001110010000:
        _o_sv = 15'b110100011100000;
      13'b1001110010001:
        _o_sv = 15'b110100011100011;
      13'b1001110010010:
        _o_sv = 15'b110100011100111;
      13'b1001110010011:
        _o_sv = 15'b110100011101011;
      13'b1001110010100:
        _o_sv = 15'b110100011101110;
      13'b1001110010101:
        _o_sv = 15'b110100011110010;
      13'b1001110010110:
        _o_sv = 15'b110100011110101;
      13'b1001110010111:
        _o_sv = 15'b110100011111001;
      13'b1001110011000:
        _o_sv = 15'b110100011111101;
      13'b1001110011001:
        _o_sv = 15'b110100100000000;
      13'b1001110011010:
        _o_sv = 15'b110100100000100;
      13'b1001110011011:
        _o_sv = 15'b110100100000111;
      13'b1001110011100:
        _o_sv = 15'b110100100001011;
      13'b1001110011101:
        _o_sv = 15'b110100100001111;
      13'b1001110011110:
        _o_sv = 15'b110100100010010;
      13'b1001110011111:
        _o_sv = 15'b110100100010110;
      13'b1001110100000:
        _o_sv = 15'b110100100011001;
      13'b1001110100001:
        _o_sv = 15'b110100100011101;
      13'b1001110100010:
        _o_sv = 15'b110100100100001;
      13'b1001110100011:
        _o_sv = 15'b110100100100100;
      13'b1001110100100:
        _o_sv = 15'b110100100101000;
      13'b1001110100101:
        _o_sv = 15'b110100100101011;
      13'b1001110100110:
        _o_sv = 15'b110100100101111;
      13'b1001110100111:
        _o_sv = 15'b110100100110010;
      13'b1001110101000:
        _o_sv = 15'b110100100110110;
      13'b1001110101001:
        _o_sv = 15'b110100100111010;
      13'b1001110101010:
        _o_sv = 15'b110100100111101;
      13'b1001110101011:
        _o_sv = 15'b110100101000001;
      13'b1001110101100:
        _o_sv = 15'b110100101000100;
      13'b1001110101101:
        _o_sv = 15'b110100101001000;
      13'b1001110101110:
        _o_sv = 15'b110100101001011;
      13'b1001110101111:
        _o_sv = 15'b110100101001111;
      13'b1001110110000:
        _o_sv = 15'b110100101010011;
      13'b1001110110001:
        _o_sv = 15'b110100101010110;
      13'b1001110110010:
        _o_sv = 15'b110100101011010;
      13'b1001110110011:
        _o_sv = 15'b110100101011101;
      13'b1001110110100:
        _o_sv = 15'b110100101100001;
      13'b1001110110101:
        _o_sv = 15'b110100101100100;
      13'b1001110110110:
        _o_sv = 15'b110100101101000;
      13'b1001110110111:
        _o_sv = 15'b110100101101100;
      13'b1001110111000:
        _o_sv = 15'b110100101101111;
      13'b1001110111001:
        _o_sv = 15'b110100101110011;
      13'b1001110111010:
        _o_sv = 15'b110100101110110;
      13'b1001110111011:
        _o_sv = 15'b110100101111010;
      13'b1001110111100:
        _o_sv = 15'b110100101111101;
      13'b1001110111101:
        _o_sv = 15'b110100110000001;
      13'b1001110111110:
        _o_sv = 15'b110100110000101;
      13'b1001110111111:
        _o_sv = 15'b110100110001000;
      13'b1001111000000:
        _o_sv = 15'b110100110001100;
      13'b1001111000001:
        _o_sv = 15'b110100110001111;
      13'b1001111000010:
        _o_sv = 15'b110100110010011;
      13'b1001111000011:
        _o_sv = 15'b110100110010110;
      13'b1001111000100:
        _o_sv = 15'b110100110011010;
      13'b1001111000101:
        _o_sv = 15'b110100110011101;
      13'b1001111000110:
        _o_sv = 15'b110100110100001;
      13'b1001111000111:
        _o_sv = 15'b110100110100101;
      13'b1001111001000:
        _o_sv = 15'b110100110101000;
      13'b1001111001001:
        _o_sv = 15'b110100110101100;
      13'b1001111001010:
        _o_sv = 15'b110100110101111;
      13'b1001111001011:
        _o_sv = 15'b110100110110011;
      13'b1001111001100:
        _o_sv = 15'b110100110110110;
      13'b1001111001101:
        _o_sv = 15'b110100110111010;
      13'b1001111001110:
        _o_sv = 15'b110100110111101;
      13'b1001111001111:
        _o_sv = 15'b110100111000001;
      13'b1001111010000:
        _o_sv = 15'b110100111000100;
      13'b1001111010001:
        _o_sv = 15'b110100111001000;
      13'b1001111010010:
        _o_sv = 15'b110100111001011;
      13'b1001111010011:
        _o_sv = 15'b110100111001111;
      13'b1001111010100:
        _o_sv = 15'b110100111010011;
      13'b1001111010101:
        _o_sv = 15'b110100111010110;
      13'b1001111010110:
        _o_sv = 15'b110100111011010;
      13'b1001111010111:
        _o_sv = 15'b110100111011101;
      13'b1001111011000:
        _o_sv = 15'b110100111100001;
      13'b1001111011001:
        _o_sv = 15'b110100111100100;
      13'b1001111011010:
        _o_sv = 15'b110100111101000;
      13'b1001111011011:
        _o_sv = 15'b110100111101011;
      13'b1001111011100:
        _o_sv = 15'b110100111101111;
      13'b1001111011101:
        _o_sv = 15'b110100111110010;
      13'b1001111011110:
        _o_sv = 15'b110100111110110;
      13'b1001111011111:
        _o_sv = 15'b110100111111001;
      13'b1001111100000:
        _o_sv = 15'b110100111111101;
      13'b1001111100001:
        _o_sv = 15'b110101000000000;
      13'b1001111100010:
        _o_sv = 15'b110101000000100;
      13'b1001111100011:
        _o_sv = 15'b110101000000111;
      13'b1001111100100:
        _o_sv = 15'b110101000001011;
      13'b1001111100101:
        _o_sv = 15'b110101000001110;
      13'b1001111100110:
        _o_sv = 15'b110101000010010;
      13'b1001111100111:
        _o_sv = 15'b110101000010110;
      13'b1001111101000:
        _o_sv = 15'b110101000011001;
      13'b1001111101001:
        _o_sv = 15'b110101000011101;
      13'b1001111101010:
        _o_sv = 15'b110101000100000;
      13'b1001111101011:
        _o_sv = 15'b110101000100100;
      13'b1001111101100:
        _o_sv = 15'b110101000100111;
      13'b1001111101101:
        _o_sv = 15'b110101000101011;
      13'b1001111101110:
        _o_sv = 15'b110101000101110;
      13'b1001111101111:
        _o_sv = 15'b110101000110010;
      13'b1001111110000:
        _o_sv = 15'b110101000110101;
      13'b1001111110001:
        _o_sv = 15'b110101000111001;
      13'b1001111110010:
        _o_sv = 15'b110101000111100;
      13'b1001111110011:
        _o_sv = 15'b110101001000000;
      13'b1001111110100:
        _o_sv = 15'b110101001000011;
      13'b1001111110101:
        _o_sv = 15'b110101001000111;
      13'b1001111110110:
        _o_sv = 15'b110101001001010;
      13'b1001111110111:
        _o_sv = 15'b110101001001110;
      13'b1001111111000:
        _o_sv = 15'b110101001010001;
      13'b1001111111001:
        _o_sv = 15'b110101001010101;
      13'b1001111111010:
        _o_sv = 15'b110101001011000;
      13'b1001111111011:
        _o_sv = 15'b110101001011100;
      13'b1001111111100:
        _o_sv = 15'b110101001011111;
      13'b1001111111101:
        _o_sv = 15'b110101001100011;
      13'b1001111111110:
        _o_sv = 15'b110101001100110;
      13'b1001111111111:
        _o_sv = 15'b110101001101010;
      13'b1010000000000:
        _o_sv = 15'b110101001101101;
      13'b1010000000001:
        _o_sv = 15'b110101001110001;
      13'b1010000000010:
        _o_sv = 15'b110101001110100;
      13'b1010000000011:
        _o_sv = 15'b110101001111000;
      13'b1010000000100:
        _o_sv = 15'b110101001111011;
      13'b1010000000101:
        _o_sv = 15'b110101001111111;
      13'b1010000000110:
        _o_sv = 15'b110101010000010;
      13'b1010000000111:
        _o_sv = 15'b110101010000110;
      13'b1010000001000:
        _o_sv = 15'b110101010001001;
      13'b1010000001001:
        _o_sv = 15'b110101010001100;
      13'b1010000001010:
        _o_sv = 15'b110101010010000;
      13'b1010000001011:
        _o_sv = 15'b110101010010011;
      13'b1010000001100:
        _o_sv = 15'b110101010010111;
      13'b1010000001101:
        _o_sv = 15'b110101010011010;
      13'b1010000001110:
        _o_sv = 15'b110101010011110;
      13'b1010000001111:
        _o_sv = 15'b110101010100001;
      13'b1010000010000:
        _o_sv = 15'b110101010100101;
      13'b1010000010001:
        _o_sv = 15'b110101010101000;
      13'b1010000010010:
        _o_sv = 15'b110101010101100;
      13'b1010000010011:
        _o_sv = 15'b110101010101111;
      13'b1010000010100:
        _o_sv = 15'b110101010110011;
      13'b1010000010101:
        _o_sv = 15'b110101010110110;
      13'b1010000010110:
        _o_sv = 15'b110101010111010;
      13'b1010000010111:
        _o_sv = 15'b110101010111101;
      13'b1010000011000:
        _o_sv = 15'b110101011000001;
      13'b1010000011001:
        _o_sv = 15'b110101011000100;
      13'b1010000011010:
        _o_sv = 15'b110101011001000;
      13'b1010000011011:
        _o_sv = 15'b110101011001011;
      13'b1010000011100:
        _o_sv = 15'b110101011001110;
      13'b1010000011101:
        _o_sv = 15'b110101011010010;
      13'b1010000011110:
        _o_sv = 15'b110101011010101;
      13'b1010000011111:
        _o_sv = 15'b110101011011001;
      13'b1010000100000:
        _o_sv = 15'b110101011011100;
      13'b1010000100001:
        _o_sv = 15'b110101011100000;
      13'b1010000100010:
        _o_sv = 15'b110101011100011;
      13'b1010000100011:
        _o_sv = 15'b110101011100111;
      13'b1010000100100:
        _o_sv = 15'b110101011101010;
      13'b1010000100101:
        _o_sv = 15'b110101011101110;
      13'b1010000100110:
        _o_sv = 15'b110101011110001;
      13'b1010000100111:
        _o_sv = 15'b110101011110100;
      13'b1010000101000:
        _o_sv = 15'b110101011111000;
      13'b1010000101001:
        _o_sv = 15'b110101011111011;
      13'b1010000101010:
        _o_sv = 15'b110101011111111;
      13'b1010000101011:
        _o_sv = 15'b110101100000010;
      13'b1010000101100:
        _o_sv = 15'b110101100000110;
      13'b1010000101101:
        _o_sv = 15'b110101100001001;
      13'b1010000101110:
        _o_sv = 15'b110101100001101;
      13'b1010000101111:
        _o_sv = 15'b110101100010000;
      13'b1010000110000:
        _o_sv = 15'b110101100010011;
      13'b1010000110001:
        _o_sv = 15'b110101100010111;
      13'b1010000110010:
        _o_sv = 15'b110101100011010;
      13'b1010000110011:
        _o_sv = 15'b110101100011110;
      13'b1010000110100:
        _o_sv = 15'b110101100100001;
      13'b1010000110101:
        _o_sv = 15'b110101100100101;
      13'b1010000110110:
        _o_sv = 15'b110101100101000;
      13'b1010000110111:
        _o_sv = 15'b110101100101100;
      13'b1010000111000:
        _o_sv = 15'b110101100101111;
      13'b1010000111001:
        _o_sv = 15'b110101100110010;
      13'b1010000111010:
        _o_sv = 15'b110101100110110;
      13'b1010000111011:
        _o_sv = 15'b110101100111001;
      13'b1010000111100:
        _o_sv = 15'b110101100111101;
      13'b1010000111101:
        _o_sv = 15'b110101101000000;
      13'b1010000111110:
        _o_sv = 15'b110101101000100;
      13'b1010000111111:
        _o_sv = 15'b110101101000111;
      13'b1010001000000:
        _o_sv = 15'b110101101001010;
      13'b1010001000001:
        _o_sv = 15'b110101101001110;
      13'b1010001000010:
        _o_sv = 15'b110101101010001;
      13'b1010001000011:
        _o_sv = 15'b110101101010101;
      13'b1010001000100:
        _o_sv = 15'b110101101011000;
      13'b1010001000101:
        _o_sv = 15'b110101101011100;
      13'b1010001000110:
        _o_sv = 15'b110101101011111;
      13'b1010001000111:
        _o_sv = 15'b110101101100010;
      13'b1010001001000:
        _o_sv = 15'b110101101100110;
      13'b1010001001001:
        _o_sv = 15'b110101101101001;
      13'b1010001001010:
        _o_sv = 15'b110101101101101;
      13'b1010001001011:
        _o_sv = 15'b110101101110000;
      13'b1010001001100:
        _o_sv = 15'b110101101110011;
      13'b1010001001101:
        _o_sv = 15'b110101101110111;
      13'b1010001001110:
        _o_sv = 15'b110101101111010;
      13'b1010001001111:
        _o_sv = 15'b110101101111110;
      13'b1010001010000:
        _o_sv = 15'b110101110000001;
      13'b1010001010001:
        _o_sv = 15'b110101110000101;
      13'b1010001010010:
        _o_sv = 15'b110101110001000;
      13'b1010001010011:
        _o_sv = 15'b110101110001011;
      13'b1010001010100:
        _o_sv = 15'b110101110001111;
      13'b1010001010101:
        _o_sv = 15'b110101110010010;
      13'b1010001010110:
        _o_sv = 15'b110101110010110;
      13'b1010001010111:
        _o_sv = 15'b110101110011001;
      13'b1010001011000:
        _o_sv = 15'b110101110011100;
      13'b1010001011001:
        _o_sv = 15'b110101110100000;
      13'b1010001011010:
        _o_sv = 15'b110101110100011;
      13'b1010001011011:
        _o_sv = 15'b110101110100111;
      13'b1010001011100:
        _o_sv = 15'b110101110101010;
      13'b1010001011101:
        _o_sv = 15'b110101110101101;
      13'b1010001011110:
        _o_sv = 15'b110101110110001;
      13'b1010001011111:
        _o_sv = 15'b110101110110100;
      13'b1010001100000:
        _o_sv = 15'b110101110111000;
      13'b1010001100001:
        _o_sv = 15'b110101110111011;
      13'b1010001100010:
        _o_sv = 15'b110101110111110;
      13'b1010001100011:
        _o_sv = 15'b110101111000010;
      13'b1010001100100:
        _o_sv = 15'b110101111000101;
      13'b1010001100101:
        _o_sv = 15'b110101111001001;
      13'b1010001100110:
        _o_sv = 15'b110101111001100;
      13'b1010001100111:
        _o_sv = 15'b110101111001111;
      13'b1010001101000:
        _o_sv = 15'b110101111010011;
      13'b1010001101001:
        _o_sv = 15'b110101111010110;
      13'b1010001101010:
        _o_sv = 15'b110101111011001;
      13'b1010001101011:
        _o_sv = 15'b110101111011101;
      13'b1010001101100:
        _o_sv = 15'b110101111100000;
      13'b1010001101101:
        _o_sv = 15'b110101111100100;
      13'b1010001101110:
        _o_sv = 15'b110101111100111;
      13'b1010001101111:
        _o_sv = 15'b110101111101010;
      13'b1010001110000:
        _o_sv = 15'b110101111101110;
      13'b1010001110001:
        _o_sv = 15'b110101111110001;
      13'b1010001110010:
        _o_sv = 15'b110101111110101;
      13'b1010001110011:
        _o_sv = 15'b110101111111000;
      13'b1010001110100:
        _o_sv = 15'b110101111111011;
      13'b1010001110101:
        _o_sv = 15'b110101111111111;
      13'b1010001110110:
        _o_sv = 15'b110110000000010;
      13'b1010001110111:
        _o_sv = 15'b110110000000101;
      13'b1010001111000:
        _o_sv = 15'b110110000001001;
      13'b1010001111001:
        _o_sv = 15'b110110000001100;
      13'b1010001111010:
        _o_sv = 15'b110110000001111;
      13'b1010001111011:
        _o_sv = 15'b110110000010011;
      13'b1010001111100:
        _o_sv = 15'b110110000010110;
      13'b1010001111101:
        _o_sv = 15'b110110000011010;
      13'b1010001111110:
        _o_sv = 15'b110110000011101;
      13'b1010001111111:
        _o_sv = 15'b110110000100000;
      13'b1010010000000:
        _o_sv = 15'b110110000100100;
      13'b1010010000001:
        _o_sv = 15'b110110000100111;
      13'b1010010000010:
        _o_sv = 15'b110110000101010;
      13'b1010010000011:
        _o_sv = 15'b110110000101110;
      13'b1010010000100:
        _o_sv = 15'b110110000110001;
      13'b1010010000101:
        _o_sv = 15'b110110000110100;
      13'b1010010000110:
        _o_sv = 15'b110110000111000;
      13'b1010010000111:
        _o_sv = 15'b110110000111011;
      13'b1010010001000:
        _o_sv = 15'b110110000111111;
      13'b1010010001001:
        _o_sv = 15'b110110001000010;
      13'b1010010001010:
        _o_sv = 15'b110110001000101;
      13'b1010010001011:
        _o_sv = 15'b110110001001001;
      13'b1010010001100:
        _o_sv = 15'b110110001001100;
      13'b1010010001101:
        _o_sv = 15'b110110001001111;
      13'b1010010001110:
        _o_sv = 15'b110110001010011;
      13'b1010010001111:
        _o_sv = 15'b110110001010110;
      13'b1010010010000:
        _o_sv = 15'b110110001011001;
      13'b1010010010001:
        _o_sv = 15'b110110001011101;
      13'b1010010010010:
        _o_sv = 15'b110110001100000;
      13'b1010010010011:
        _o_sv = 15'b110110001100011;
      13'b1010010010100:
        _o_sv = 15'b110110001100111;
      13'b1010010010101:
        _o_sv = 15'b110110001101010;
      13'b1010010010110:
        _o_sv = 15'b110110001101101;
      13'b1010010010111:
        _o_sv = 15'b110110001110001;
      13'b1010010011000:
        _o_sv = 15'b110110001110100;
      13'b1010010011001:
        _o_sv = 15'b110110001110111;
      13'b1010010011010:
        _o_sv = 15'b110110001111011;
      13'b1010010011011:
        _o_sv = 15'b110110001111110;
      13'b1010010011100:
        _o_sv = 15'b110110010000001;
      13'b1010010011101:
        _o_sv = 15'b110110010000101;
      13'b1010010011110:
        _o_sv = 15'b110110010001000;
      13'b1010010011111:
        _o_sv = 15'b110110010001011;
      13'b1010010100000:
        _o_sv = 15'b110110010001111;
      13'b1010010100001:
        _o_sv = 15'b110110010010010;
      13'b1010010100010:
        _o_sv = 15'b110110010010101;
      13'b1010010100011:
        _o_sv = 15'b110110010011001;
      13'b1010010100100:
        _o_sv = 15'b110110010011100;
      13'b1010010100101:
        _o_sv = 15'b110110010011111;
      13'b1010010100110:
        _o_sv = 15'b110110010100011;
      13'b1010010100111:
        _o_sv = 15'b110110010100110;
      13'b1010010101000:
        _o_sv = 15'b110110010101001;
      13'b1010010101001:
        _o_sv = 15'b110110010101101;
      13'b1010010101010:
        _o_sv = 15'b110110010110000;
      13'b1010010101011:
        _o_sv = 15'b110110010110011;
      13'b1010010101100:
        _o_sv = 15'b110110010110111;
      13'b1010010101101:
        _o_sv = 15'b110110010111010;
      13'b1010010101110:
        _o_sv = 15'b110110010111101;
      13'b1010010101111:
        _o_sv = 15'b110110011000001;
      13'b1010010110000:
        _o_sv = 15'b110110011000100;
      13'b1010010110001:
        _o_sv = 15'b110110011000111;
      13'b1010010110010:
        _o_sv = 15'b110110011001010;
      13'b1010010110011:
        _o_sv = 15'b110110011001110;
      13'b1010010110100:
        _o_sv = 15'b110110011010001;
      13'b1010010110101:
        _o_sv = 15'b110110011010100;
      13'b1010010110110:
        _o_sv = 15'b110110011011000;
      13'b1010010110111:
        _o_sv = 15'b110110011011011;
      13'b1010010111000:
        _o_sv = 15'b110110011011110;
      13'b1010010111001:
        _o_sv = 15'b110110011100010;
      13'b1010010111010:
        _o_sv = 15'b110110011100101;
      13'b1010010111011:
        _o_sv = 15'b110110011101000;
      13'b1010010111100:
        _o_sv = 15'b110110011101100;
      13'b1010010111101:
        _o_sv = 15'b110110011101111;
      13'b1010010111110:
        _o_sv = 15'b110110011110010;
      13'b1010010111111:
        _o_sv = 15'b110110011110101;
      13'b1010011000000:
        _o_sv = 15'b110110011111001;
      13'b1010011000001:
        _o_sv = 15'b110110011111100;
      13'b1010011000010:
        _o_sv = 15'b110110011111111;
      13'b1010011000011:
        _o_sv = 15'b110110100000011;
      13'b1010011000100:
        _o_sv = 15'b110110100000110;
      13'b1010011000101:
        _o_sv = 15'b110110100001001;
      13'b1010011000110:
        _o_sv = 15'b110110100001100;
      13'b1010011000111:
        _o_sv = 15'b110110100010000;
      13'b1010011001000:
        _o_sv = 15'b110110100010011;
      13'b1010011001001:
        _o_sv = 15'b110110100010110;
      13'b1010011001010:
        _o_sv = 15'b110110100011010;
      13'b1010011001011:
        _o_sv = 15'b110110100011101;
      13'b1010011001100:
        _o_sv = 15'b110110100100000;
      13'b1010011001101:
        _o_sv = 15'b110110100100011;
      13'b1010011001110:
        _o_sv = 15'b110110100100111;
      13'b1010011001111:
        _o_sv = 15'b110110100101010;
      13'b1010011010000:
        _o_sv = 15'b110110100101101;
      13'b1010011010001:
        _o_sv = 15'b110110100110001;
      13'b1010011010010:
        _o_sv = 15'b110110100110100;
      13'b1010011010011:
        _o_sv = 15'b110110100110111;
      13'b1010011010100:
        _o_sv = 15'b110110100111010;
      13'b1010011010101:
        _o_sv = 15'b110110100111110;
      13'b1010011010110:
        _o_sv = 15'b110110101000001;
      13'b1010011010111:
        _o_sv = 15'b110110101000100;
      13'b1010011011000:
        _o_sv = 15'b110110101001000;
      13'b1010011011001:
        _o_sv = 15'b110110101001011;
      13'b1010011011010:
        _o_sv = 15'b110110101001110;
      13'b1010011011011:
        _o_sv = 15'b110110101010001;
      13'b1010011011100:
        _o_sv = 15'b110110101010101;
      13'b1010011011101:
        _o_sv = 15'b110110101011000;
      13'b1010011011110:
        _o_sv = 15'b110110101011011;
      13'b1010011011111:
        _o_sv = 15'b110110101011110;
      13'b1010011100000:
        _o_sv = 15'b110110101100010;
      13'b1010011100001:
        _o_sv = 15'b110110101100101;
      13'b1010011100010:
        _o_sv = 15'b110110101101000;
      13'b1010011100011:
        _o_sv = 15'b110110101101011;
      13'b1010011100100:
        _o_sv = 15'b110110101101111;
      13'b1010011100101:
        _o_sv = 15'b110110101110010;
      13'b1010011100110:
        _o_sv = 15'b110110101110101;
      13'b1010011100111:
        _o_sv = 15'b110110101111000;
      13'b1010011101000:
        _o_sv = 15'b110110101111100;
      13'b1010011101001:
        _o_sv = 15'b110110101111111;
      13'b1010011101010:
        _o_sv = 15'b110110110000010;
      13'b1010011101011:
        _o_sv = 15'b110110110000101;
      13'b1010011101100:
        _o_sv = 15'b110110110001001;
      13'b1010011101101:
        _o_sv = 15'b110110110001100;
      13'b1010011101110:
        _o_sv = 15'b110110110001111;
      13'b1010011101111:
        _o_sv = 15'b110110110010010;
      13'b1010011110000:
        _o_sv = 15'b110110110010110;
      13'b1010011110001:
        _o_sv = 15'b110110110011001;
      13'b1010011110010:
        _o_sv = 15'b110110110011100;
      13'b1010011110011:
        _o_sv = 15'b110110110011111;
      13'b1010011110100:
        _o_sv = 15'b110110110100011;
      13'b1010011110101:
        _o_sv = 15'b110110110100110;
      13'b1010011110110:
        _o_sv = 15'b110110110101001;
      13'b1010011110111:
        _o_sv = 15'b110110110101100;
      13'b1010011111000:
        _o_sv = 15'b110110110110000;
      13'b1010011111001:
        _o_sv = 15'b110110110110011;
      13'b1010011111010:
        _o_sv = 15'b110110110110110;
      13'b1010011111011:
        _o_sv = 15'b110110110111001;
      13'b1010011111100:
        _o_sv = 15'b110110110111101;
      13'b1010011111101:
        _o_sv = 15'b110110111000000;
      13'b1010011111110:
        _o_sv = 15'b110110111000011;
      13'b1010011111111:
        _o_sv = 15'b110110111000110;
      13'b1010100000000:
        _o_sv = 15'b110110111001010;
      13'b1010100000001:
        _o_sv = 15'b110110111001101;
      13'b1010100000010:
        _o_sv = 15'b110110111010000;
      13'b1010100000011:
        _o_sv = 15'b110110111010011;
      13'b1010100000100:
        _o_sv = 15'b110110111010110;
      13'b1010100000101:
        _o_sv = 15'b110110111011010;
      13'b1010100000110:
        _o_sv = 15'b110110111011101;
      13'b1010100000111:
        _o_sv = 15'b110110111100000;
      13'b1010100001000:
        _o_sv = 15'b110110111100011;
      13'b1010100001001:
        _o_sv = 15'b110110111100111;
      13'b1010100001010:
        _o_sv = 15'b110110111101010;
      13'b1010100001011:
        _o_sv = 15'b110110111101101;
      13'b1010100001100:
        _o_sv = 15'b110110111110000;
      13'b1010100001101:
        _o_sv = 15'b110110111110011;
      13'b1010100001110:
        _o_sv = 15'b110110111110111;
      13'b1010100001111:
        _o_sv = 15'b110110111111010;
      13'b1010100010000:
        _o_sv = 15'b110110111111101;
      13'b1010100010001:
        _o_sv = 15'b110111000000000;
      13'b1010100010010:
        _o_sv = 15'b110111000000100;
      13'b1010100010011:
        _o_sv = 15'b110111000000111;
      13'b1010100010100:
        _o_sv = 15'b110111000001010;
      13'b1010100010101:
        _o_sv = 15'b110111000001101;
      13'b1010100010110:
        _o_sv = 15'b110111000010000;
      13'b1010100010111:
        _o_sv = 15'b110111000010100;
      13'b1010100011000:
        _o_sv = 15'b110111000010111;
      13'b1010100011001:
        _o_sv = 15'b110111000011010;
      13'b1010100011010:
        _o_sv = 15'b110111000011101;
      13'b1010100011011:
        _o_sv = 15'b110111000100000;
      13'b1010100011100:
        _o_sv = 15'b110111000100100;
      13'b1010100011101:
        _o_sv = 15'b110111000100111;
      13'b1010100011110:
        _o_sv = 15'b110111000101010;
      13'b1010100011111:
        _o_sv = 15'b110111000101101;
      13'b1010100100000:
        _o_sv = 15'b110111000110000;
      13'b1010100100001:
        _o_sv = 15'b110111000110100;
      13'b1010100100010:
        _o_sv = 15'b110111000110111;
      13'b1010100100011:
        _o_sv = 15'b110111000111010;
      13'b1010100100100:
        _o_sv = 15'b110111000111101;
      13'b1010100100101:
        _o_sv = 15'b110111001000000;
      13'b1010100100110:
        _o_sv = 15'b110111001000100;
      13'b1010100100111:
        _o_sv = 15'b110111001000111;
      13'b1010100101000:
        _o_sv = 15'b110111001001010;
      13'b1010100101001:
        _o_sv = 15'b110111001001101;
      13'b1010100101010:
        _o_sv = 15'b110111001010000;
      13'b1010100101011:
        _o_sv = 15'b110111001010011;
      13'b1010100101100:
        _o_sv = 15'b110111001010111;
      13'b1010100101101:
        _o_sv = 15'b110111001011010;
      13'b1010100101110:
        _o_sv = 15'b110111001011101;
      13'b1010100101111:
        _o_sv = 15'b110111001100000;
      13'b1010100110000:
        _o_sv = 15'b110111001100011;
      13'b1010100110001:
        _o_sv = 15'b110111001100111;
      13'b1010100110010:
        _o_sv = 15'b110111001101010;
      13'b1010100110011:
        _o_sv = 15'b110111001101101;
      13'b1010100110100:
        _o_sv = 15'b110111001110000;
      13'b1010100110101:
        _o_sv = 15'b110111001110011;
      13'b1010100110110:
        _o_sv = 15'b110111001110110;
      13'b1010100110111:
        _o_sv = 15'b110111001111010;
      13'b1010100111000:
        _o_sv = 15'b110111001111101;
      13'b1010100111001:
        _o_sv = 15'b110111010000000;
      13'b1010100111010:
        _o_sv = 15'b110111010000011;
      13'b1010100111011:
        _o_sv = 15'b110111010000110;
      13'b1010100111100:
        _o_sv = 15'b110111010001001;
      13'b1010100111101:
        _o_sv = 15'b110111010001101;
      13'b1010100111110:
        _o_sv = 15'b110111010010000;
      13'b1010100111111:
        _o_sv = 15'b110111010010011;
      13'b1010101000000:
        _o_sv = 15'b110111010010110;
      13'b1010101000001:
        _o_sv = 15'b110111010011001;
      13'b1010101000010:
        _o_sv = 15'b110111010011100;
      13'b1010101000011:
        _o_sv = 15'b110111010100000;
      13'b1010101000100:
        _o_sv = 15'b110111010100011;
      13'b1010101000101:
        _o_sv = 15'b110111010100110;
      13'b1010101000110:
        _o_sv = 15'b110111010101001;
      13'b1010101000111:
        _o_sv = 15'b110111010101100;
      13'b1010101001000:
        _o_sv = 15'b110111010101111;
      13'b1010101001001:
        _o_sv = 15'b110111010110011;
      13'b1010101001010:
        _o_sv = 15'b110111010110110;
      13'b1010101001011:
        _o_sv = 15'b110111010111001;
      13'b1010101001100:
        _o_sv = 15'b110111010111100;
      13'b1010101001101:
        _o_sv = 15'b110111010111111;
      13'b1010101001110:
        _o_sv = 15'b110111011000010;
      13'b1010101001111:
        _o_sv = 15'b110111011000110;
      13'b1010101010000:
        _o_sv = 15'b110111011001001;
      13'b1010101010001:
        _o_sv = 15'b110111011001100;
      13'b1010101010010:
        _o_sv = 15'b110111011001111;
      13'b1010101010011:
        _o_sv = 15'b110111011010010;
      13'b1010101010100:
        _o_sv = 15'b110111011010101;
      13'b1010101010101:
        _o_sv = 15'b110111011011000;
      13'b1010101010110:
        _o_sv = 15'b110111011011100;
      13'b1010101010111:
        _o_sv = 15'b110111011011111;
      13'b1010101011000:
        _o_sv = 15'b110111011100010;
      13'b1010101011001:
        _o_sv = 15'b110111011100101;
      13'b1010101011010:
        _o_sv = 15'b110111011101000;
      13'b1010101011011:
        _o_sv = 15'b110111011101011;
      13'b1010101011100:
        _o_sv = 15'b110111011101110;
      13'b1010101011101:
        _o_sv = 15'b110111011110001;
      13'b1010101011110:
        _o_sv = 15'b110111011110101;
      13'b1010101011111:
        _o_sv = 15'b110111011111000;
      13'b1010101100000:
        _o_sv = 15'b110111011111011;
      13'b1010101100001:
        _o_sv = 15'b110111011111110;
      13'b1010101100010:
        _o_sv = 15'b110111100000001;
      13'b1010101100011:
        _o_sv = 15'b110111100000100;
      13'b1010101100100:
        _o_sv = 15'b110111100000111;
      13'b1010101100101:
        _o_sv = 15'b110111100001011;
      13'b1010101100110:
        _o_sv = 15'b110111100001110;
      13'b1010101100111:
        _o_sv = 15'b110111100010001;
      13'b1010101101000:
        _o_sv = 15'b110111100010100;
      13'b1010101101001:
        _o_sv = 15'b110111100010111;
      13'b1010101101010:
        _o_sv = 15'b110111100011010;
      13'b1010101101011:
        _o_sv = 15'b110111100011101;
      13'b1010101101100:
        _o_sv = 15'b110111100100000;
      13'b1010101101101:
        _o_sv = 15'b110111100100011;
      13'b1010101101110:
        _o_sv = 15'b110111100100111;
      13'b1010101101111:
        _o_sv = 15'b110111100101010;
      13'b1010101110000:
        _o_sv = 15'b110111100101101;
      13'b1010101110001:
        _o_sv = 15'b110111100110000;
      13'b1010101110010:
        _o_sv = 15'b110111100110011;
      13'b1010101110011:
        _o_sv = 15'b110111100110110;
      13'b1010101110100:
        _o_sv = 15'b110111100111001;
      13'b1010101110101:
        _o_sv = 15'b110111100111100;
      13'b1010101110110:
        _o_sv = 15'b110111100111111;
      13'b1010101110111:
        _o_sv = 15'b110111101000011;
      13'b1010101111000:
        _o_sv = 15'b110111101000110;
      13'b1010101111001:
        _o_sv = 15'b110111101001001;
      13'b1010101111010:
        _o_sv = 15'b110111101001100;
      13'b1010101111011:
        _o_sv = 15'b110111101001111;
      13'b1010101111100:
        _o_sv = 15'b110111101010010;
      13'b1010101111101:
        _o_sv = 15'b110111101010101;
      13'b1010101111110:
        _o_sv = 15'b110111101011000;
      13'b1010101111111:
        _o_sv = 15'b110111101011011;
      13'b1010110000000:
        _o_sv = 15'b110111101011111;
      13'b1010110000001:
        _o_sv = 15'b110111101100010;
      13'b1010110000010:
        _o_sv = 15'b110111101100101;
      13'b1010110000011:
        _o_sv = 15'b110111101101000;
      13'b1010110000100:
        _o_sv = 15'b110111101101011;
      13'b1010110000101:
        _o_sv = 15'b110111101101110;
      13'b1010110000110:
        _o_sv = 15'b110111101110001;
      13'b1010110000111:
        _o_sv = 15'b110111101110100;
      13'b1010110001000:
        _o_sv = 15'b110111101110111;
      13'b1010110001001:
        _o_sv = 15'b110111101111010;
      13'b1010110001010:
        _o_sv = 15'b110111101111101;
      13'b1010110001011:
        _o_sv = 15'b110111110000001;
      13'b1010110001100:
        _o_sv = 15'b110111110000100;
      13'b1010110001101:
        _o_sv = 15'b110111110000111;
      13'b1010110001110:
        _o_sv = 15'b110111110001010;
      13'b1010110001111:
        _o_sv = 15'b110111110001101;
      13'b1010110010000:
        _o_sv = 15'b110111110010000;
      13'b1010110010001:
        _o_sv = 15'b110111110010011;
      13'b1010110010010:
        _o_sv = 15'b110111110010110;
      13'b1010110010011:
        _o_sv = 15'b110111110011001;
      13'b1010110010100:
        _o_sv = 15'b110111110011100;
      13'b1010110010101:
        _o_sv = 15'b110111110011111;
      13'b1010110010110:
        _o_sv = 15'b110111110100010;
      13'b1010110010111:
        _o_sv = 15'b110111110100101;
      13'b1010110011000:
        _o_sv = 15'b110111110101001;
      13'b1010110011001:
        _o_sv = 15'b110111110101100;
      13'b1010110011010:
        _o_sv = 15'b110111110101111;
      13'b1010110011011:
        _o_sv = 15'b110111110110010;
      13'b1010110011100:
        _o_sv = 15'b110111110110101;
      13'b1010110011101:
        _o_sv = 15'b110111110111000;
      13'b1010110011110:
        _o_sv = 15'b110111110111011;
      13'b1010110011111:
        _o_sv = 15'b110111110111110;
      13'b1010110100000:
        _o_sv = 15'b110111111000001;
      13'b1010110100001:
        _o_sv = 15'b110111111000100;
      13'b1010110100010:
        _o_sv = 15'b110111111000111;
      13'b1010110100011:
        _o_sv = 15'b110111111001010;
      13'b1010110100100:
        _o_sv = 15'b110111111001101;
      13'b1010110100101:
        _o_sv = 15'b110111111010000;
      13'b1010110100110:
        _o_sv = 15'b110111111010011;
      13'b1010110100111:
        _o_sv = 15'b110111111010110;
      13'b1010110101000:
        _o_sv = 15'b110111111011010;
      13'b1010110101001:
        _o_sv = 15'b110111111011101;
      13'b1010110101010:
        _o_sv = 15'b110111111100000;
      13'b1010110101011:
        _o_sv = 15'b110111111100011;
      13'b1010110101100:
        _o_sv = 15'b110111111100110;
      13'b1010110101101:
        _o_sv = 15'b110111111101001;
      13'b1010110101110:
        _o_sv = 15'b110111111101100;
      13'b1010110101111:
        _o_sv = 15'b110111111101111;
      13'b1010110110000:
        _o_sv = 15'b110111111110010;
      13'b1010110110001:
        _o_sv = 15'b110111111110101;
      13'b1010110110010:
        _o_sv = 15'b110111111111000;
      13'b1010110110011:
        _o_sv = 15'b110111111111011;
      13'b1010110110100:
        _o_sv = 15'b110111111111110;
      13'b1010110110101:
        _o_sv = 15'b111000000000001;
      13'b1010110110110:
        _o_sv = 15'b111000000000100;
      13'b1010110110111:
        _o_sv = 15'b111000000000111;
      13'b1010110111000:
        _o_sv = 15'b111000000001010;
      13'b1010110111001:
        _o_sv = 15'b111000000001101;
      13'b1010110111010:
        _o_sv = 15'b111000000010000;
      13'b1010110111011:
        _o_sv = 15'b111000000010011;
      13'b1010110111100:
        _o_sv = 15'b111000000010110;
      13'b1010110111101:
        _o_sv = 15'b111000000011001;
      13'b1010110111110:
        _o_sv = 15'b111000000011101;
      13'b1010110111111:
        _o_sv = 15'b111000000100000;
      13'b1010111000000:
        _o_sv = 15'b111000000100011;
      13'b1010111000001:
        _o_sv = 15'b111000000100110;
      13'b1010111000010:
        _o_sv = 15'b111000000101001;
      13'b1010111000011:
        _o_sv = 15'b111000000101100;
      13'b1010111000100:
        _o_sv = 15'b111000000101111;
      13'b1010111000101:
        _o_sv = 15'b111000000110010;
      13'b1010111000110:
        _o_sv = 15'b111000000110101;
      13'b1010111000111:
        _o_sv = 15'b111000000111000;
      13'b1010111001000:
        _o_sv = 15'b111000000111011;
      13'b1010111001001:
        _o_sv = 15'b111000000111110;
      13'b1010111001010:
        _o_sv = 15'b111000001000001;
      13'b1010111001011:
        _o_sv = 15'b111000001000100;
      13'b1010111001100:
        _o_sv = 15'b111000001000111;
      13'b1010111001101:
        _o_sv = 15'b111000001001010;
      13'b1010111001110:
        _o_sv = 15'b111000001001101;
      13'b1010111001111:
        _o_sv = 15'b111000001010000;
      13'b1010111010000:
        _o_sv = 15'b111000001010011;
      13'b1010111010001:
        _o_sv = 15'b111000001010110;
      13'b1010111010010:
        _o_sv = 15'b111000001011001;
      13'b1010111010011:
        _o_sv = 15'b111000001011100;
      13'b1010111010100:
        _o_sv = 15'b111000001011111;
      13'b1010111010101:
        _o_sv = 15'b111000001100010;
      13'b1010111010110:
        _o_sv = 15'b111000001100101;
      13'b1010111010111:
        _o_sv = 15'b111000001101000;
      13'b1010111011000:
        _o_sv = 15'b111000001101011;
      13'b1010111011001:
        _o_sv = 15'b111000001101110;
      13'b1010111011010:
        _o_sv = 15'b111000001110001;
      13'b1010111011011:
        _o_sv = 15'b111000001110100;
      13'b1010111011100:
        _o_sv = 15'b111000001110111;
      13'b1010111011101:
        _o_sv = 15'b111000001111010;
      13'b1010111011110:
        _o_sv = 15'b111000001111101;
      13'b1010111011111:
        _o_sv = 15'b111000010000000;
      13'b1010111100000:
        _o_sv = 15'b111000010000011;
      13'b1010111100001:
        _o_sv = 15'b111000010000110;
      13'b1010111100010:
        _o_sv = 15'b111000010001001;
      13'b1010111100011:
        _o_sv = 15'b111000010001100;
      13'b1010111100100:
        _o_sv = 15'b111000010001111;
      13'b1010111100101:
        _o_sv = 15'b111000010010010;
      13'b1010111100110:
        _o_sv = 15'b111000010010101;
      13'b1010111100111:
        _o_sv = 15'b111000010011000;
      13'b1010111101000:
        _o_sv = 15'b111000010011011;
      13'b1010111101001:
        _o_sv = 15'b111000010011110;
      13'b1010111101010:
        _o_sv = 15'b111000010100001;
      13'b1010111101011:
        _o_sv = 15'b111000010100100;
      13'b1010111101100:
        _o_sv = 15'b111000010100111;
      13'b1010111101101:
        _o_sv = 15'b111000010101010;
      13'b1010111101110:
        _o_sv = 15'b111000010101101;
      13'b1010111101111:
        _o_sv = 15'b111000010110000;
      13'b1010111110000:
        _o_sv = 15'b111000010110011;
      13'b1010111110001:
        _o_sv = 15'b111000010110110;
      13'b1010111110010:
        _o_sv = 15'b111000010111001;
      13'b1010111110011:
        _o_sv = 15'b111000010111100;
      13'b1010111110100:
        _o_sv = 15'b111000010111111;
      13'b1010111110101:
        _o_sv = 15'b111000011000010;
      13'b1010111110110:
        _o_sv = 15'b111000011000101;
      13'b1010111110111:
        _o_sv = 15'b111000011001000;
      13'b1010111111000:
        _o_sv = 15'b111000011001011;
      13'b1010111111001:
        _o_sv = 15'b111000011001110;
      13'b1010111111010:
        _o_sv = 15'b111000011010001;
      13'b1010111111011:
        _o_sv = 15'b111000011010011;
      13'b1010111111100:
        _o_sv = 15'b111000011010110;
      13'b1010111111101:
        _o_sv = 15'b111000011011001;
      13'b1010111111110:
        _o_sv = 15'b111000011011100;
      13'b1010111111111:
        _o_sv = 15'b111000011011111;
      13'b1011000000000:
        _o_sv = 15'b111000011100010;
      13'b1011000000001:
        _o_sv = 15'b111000011100101;
      13'b1011000000010:
        _o_sv = 15'b111000011101000;
      13'b1011000000011:
        _o_sv = 15'b111000011101011;
      13'b1011000000100:
        _o_sv = 15'b111000011101110;
      13'b1011000000101:
        _o_sv = 15'b111000011110001;
      13'b1011000000110:
        _o_sv = 15'b111000011110100;
      13'b1011000000111:
        _o_sv = 15'b111000011110111;
      13'b1011000001000:
        _o_sv = 15'b111000011111010;
      13'b1011000001001:
        _o_sv = 15'b111000011111101;
      13'b1011000001010:
        _o_sv = 15'b111000100000000;
      13'b1011000001011:
        _o_sv = 15'b111000100000011;
      13'b1011000001100:
        _o_sv = 15'b111000100000110;
      13'b1011000001101:
        _o_sv = 15'b111000100001001;
      13'b1011000001110:
        _o_sv = 15'b111000100001100;
      13'b1011000001111:
        _o_sv = 15'b111000100001111;
      13'b1011000010000:
        _o_sv = 15'b111000100010010;
      13'b1011000010001:
        _o_sv = 15'b111000100010100;
      13'b1011000010010:
        _o_sv = 15'b111000100010111;
      13'b1011000010011:
        _o_sv = 15'b111000100011010;
      13'b1011000010100:
        _o_sv = 15'b111000100011101;
      13'b1011000010101:
        _o_sv = 15'b111000100100000;
      13'b1011000010110:
        _o_sv = 15'b111000100100011;
      13'b1011000010111:
        _o_sv = 15'b111000100100110;
      13'b1011000011000:
        _o_sv = 15'b111000100101001;
      13'b1011000011001:
        _o_sv = 15'b111000100101100;
      13'b1011000011010:
        _o_sv = 15'b111000100101111;
      13'b1011000011011:
        _o_sv = 15'b111000100110010;
      13'b1011000011100:
        _o_sv = 15'b111000100110101;
      13'b1011000011101:
        _o_sv = 15'b111000100111000;
      13'b1011000011110:
        _o_sv = 15'b111000100111011;
      13'b1011000011111:
        _o_sv = 15'b111000100111110;
      13'b1011000100000:
        _o_sv = 15'b111000101000001;
      13'b1011000100001:
        _o_sv = 15'b111000101000011;
      13'b1011000100010:
        _o_sv = 15'b111000101000110;
      13'b1011000100011:
        _o_sv = 15'b111000101001001;
      13'b1011000100100:
        _o_sv = 15'b111000101001100;
      13'b1011000100101:
        _o_sv = 15'b111000101001111;
      13'b1011000100110:
        _o_sv = 15'b111000101010010;
      13'b1011000100111:
        _o_sv = 15'b111000101010101;
      13'b1011000101000:
        _o_sv = 15'b111000101011000;
      13'b1011000101001:
        _o_sv = 15'b111000101011011;
      13'b1011000101010:
        _o_sv = 15'b111000101011110;
      13'b1011000101011:
        _o_sv = 15'b111000101100001;
      13'b1011000101100:
        _o_sv = 15'b111000101100100;
      13'b1011000101101:
        _o_sv = 15'b111000101100111;
      13'b1011000101110:
        _o_sv = 15'b111000101101001;
      13'b1011000101111:
        _o_sv = 15'b111000101101100;
      13'b1011000110000:
        _o_sv = 15'b111000101101111;
      13'b1011000110001:
        _o_sv = 15'b111000101110010;
      13'b1011000110010:
        _o_sv = 15'b111000101110101;
      13'b1011000110011:
        _o_sv = 15'b111000101111000;
      13'b1011000110100:
        _o_sv = 15'b111000101111011;
      13'b1011000110101:
        _o_sv = 15'b111000101111110;
      13'b1011000110110:
        _o_sv = 15'b111000110000001;
      13'b1011000110111:
        _o_sv = 15'b111000110000100;
      13'b1011000111000:
        _o_sv = 15'b111000110000110;
      13'b1011000111001:
        _o_sv = 15'b111000110001001;
      13'b1011000111010:
        _o_sv = 15'b111000110001100;
      13'b1011000111011:
        _o_sv = 15'b111000110001111;
      13'b1011000111100:
        _o_sv = 15'b111000110010010;
      13'b1011000111101:
        _o_sv = 15'b111000110010101;
      13'b1011000111110:
        _o_sv = 15'b111000110011000;
      13'b1011000111111:
        _o_sv = 15'b111000110011011;
      13'b1011001000000:
        _o_sv = 15'b111000110011110;
      13'b1011001000001:
        _o_sv = 15'b111000110100001;
      13'b1011001000010:
        _o_sv = 15'b111000110100011;
      13'b1011001000011:
        _o_sv = 15'b111000110100110;
      13'b1011001000100:
        _o_sv = 15'b111000110101001;
      13'b1011001000101:
        _o_sv = 15'b111000110101100;
      13'b1011001000110:
        _o_sv = 15'b111000110101111;
      13'b1011001000111:
        _o_sv = 15'b111000110110010;
      13'b1011001001000:
        _o_sv = 15'b111000110110101;
      13'b1011001001001:
        _o_sv = 15'b111000110111000;
      13'b1011001001010:
        _o_sv = 15'b111000110111011;
      13'b1011001001011:
        _o_sv = 15'b111000110111101;
      13'b1011001001100:
        _o_sv = 15'b111000111000000;
      13'b1011001001101:
        _o_sv = 15'b111000111000011;
      13'b1011001001110:
        _o_sv = 15'b111000111000110;
      13'b1011001001111:
        _o_sv = 15'b111000111001001;
      13'b1011001010000:
        _o_sv = 15'b111000111001100;
      13'b1011001010001:
        _o_sv = 15'b111000111001111;
      13'b1011001010010:
        _o_sv = 15'b111000111010010;
      13'b1011001010011:
        _o_sv = 15'b111000111010100;
      13'b1011001010100:
        _o_sv = 15'b111000111010111;
      13'b1011001010101:
        _o_sv = 15'b111000111011010;
      13'b1011001010110:
        _o_sv = 15'b111000111011101;
      13'b1011001010111:
        _o_sv = 15'b111000111100000;
      13'b1011001011000:
        _o_sv = 15'b111000111100011;
      13'b1011001011001:
        _o_sv = 15'b111000111100110;
      13'b1011001011010:
        _o_sv = 15'b111000111101001;
      13'b1011001011011:
        _o_sv = 15'b111000111101011;
      13'b1011001011100:
        _o_sv = 15'b111000111101110;
      13'b1011001011101:
        _o_sv = 15'b111000111110001;
      13'b1011001011110:
        _o_sv = 15'b111000111110100;
      13'b1011001011111:
        _o_sv = 15'b111000111110111;
      13'b1011001100000:
        _o_sv = 15'b111000111111010;
      13'b1011001100001:
        _o_sv = 15'b111000111111101;
      13'b1011001100010:
        _o_sv = 15'b111000111111111;
      13'b1011001100011:
        _o_sv = 15'b111001000000010;
      13'b1011001100100:
        _o_sv = 15'b111001000000101;
      13'b1011001100101:
        _o_sv = 15'b111001000001000;
      13'b1011001100110:
        _o_sv = 15'b111001000001011;
      13'b1011001100111:
        _o_sv = 15'b111001000001110;
      13'b1011001101000:
        _o_sv = 15'b111001000010001;
      13'b1011001101001:
        _o_sv = 15'b111001000010011;
      13'b1011001101010:
        _o_sv = 15'b111001000010110;
      13'b1011001101011:
        _o_sv = 15'b111001000011001;
      13'b1011001101100:
        _o_sv = 15'b111001000011100;
      13'b1011001101101:
        _o_sv = 15'b111001000011111;
      13'b1011001101110:
        _o_sv = 15'b111001000100010;
      13'b1011001101111:
        _o_sv = 15'b111001000100100;
      13'b1011001110000:
        _o_sv = 15'b111001000100111;
      13'b1011001110001:
        _o_sv = 15'b111001000101010;
      13'b1011001110010:
        _o_sv = 15'b111001000101101;
      13'b1011001110011:
        _o_sv = 15'b111001000110000;
      13'b1011001110100:
        _o_sv = 15'b111001000110011;
      13'b1011001110101:
        _o_sv = 15'b111001000110110;
      13'b1011001110110:
        _o_sv = 15'b111001000111000;
      13'b1011001110111:
        _o_sv = 15'b111001000111011;
      13'b1011001111000:
        _o_sv = 15'b111001000111110;
      13'b1011001111001:
        _o_sv = 15'b111001001000001;
      13'b1011001111010:
        _o_sv = 15'b111001001000100;
      13'b1011001111011:
        _o_sv = 15'b111001001000111;
      13'b1011001111100:
        _o_sv = 15'b111001001001001;
      13'b1011001111101:
        _o_sv = 15'b111001001001100;
      13'b1011001111110:
        _o_sv = 15'b111001001001111;
      13'b1011001111111:
        _o_sv = 15'b111001001010010;
      13'b1011010000000:
        _o_sv = 15'b111001001010101;
      13'b1011010000001:
        _o_sv = 15'b111001001010111;
      13'b1011010000010:
        _o_sv = 15'b111001001011010;
      13'b1011010000011:
        _o_sv = 15'b111001001011101;
      13'b1011010000100:
        _o_sv = 15'b111001001100000;
      13'b1011010000101:
        _o_sv = 15'b111001001100011;
      13'b1011010000110:
        _o_sv = 15'b111001001100110;
      13'b1011010000111:
        _o_sv = 15'b111001001101000;
      13'b1011010001000:
        _o_sv = 15'b111001001101011;
      13'b1011010001001:
        _o_sv = 15'b111001001101110;
      13'b1011010001010:
        _o_sv = 15'b111001001110001;
      13'b1011010001011:
        _o_sv = 15'b111001001110100;
      13'b1011010001100:
        _o_sv = 15'b111001001110110;
      13'b1011010001101:
        _o_sv = 15'b111001001111001;
      13'b1011010001110:
        _o_sv = 15'b111001001111100;
      13'b1011010001111:
        _o_sv = 15'b111001001111111;
      13'b1011010010000:
        _o_sv = 15'b111001010000010;
      13'b1011010010001:
        _o_sv = 15'b111001010000101;
      13'b1011010010010:
        _o_sv = 15'b111001010000111;
      13'b1011010010011:
        _o_sv = 15'b111001010001010;
      13'b1011010010100:
        _o_sv = 15'b111001010001101;
      13'b1011010010101:
        _o_sv = 15'b111001010010000;
      13'b1011010010110:
        _o_sv = 15'b111001010010011;
      13'b1011010010111:
        _o_sv = 15'b111001010010101;
      13'b1011010011000:
        _o_sv = 15'b111001010011000;
      13'b1011010011001:
        _o_sv = 15'b111001010011011;
      13'b1011010011010:
        _o_sv = 15'b111001010011110;
      13'b1011010011011:
        _o_sv = 15'b111001010100001;
      13'b1011010011100:
        _o_sv = 15'b111001010100011;
      13'b1011010011101:
        _o_sv = 15'b111001010100110;
      13'b1011010011110:
        _o_sv = 15'b111001010101001;
      13'b1011010011111:
        _o_sv = 15'b111001010101100;
      13'b1011010100000:
        _o_sv = 15'b111001010101111;
      13'b1011010100001:
        _o_sv = 15'b111001010110001;
      13'b1011010100010:
        _o_sv = 15'b111001010110100;
      13'b1011010100011:
        _o_sv = 15'b111001010110111;
      13'b1011010100100:
        _o_sv = 15'b111001010111010;
      13'b1011010100101:
        _o_sv = 15'b111001010111100;
      13'b1011010100110:
        _o_sv = 15'b111001010111111;
      13'b1011010100111:
        _o_sv = 15'b111001011000010;
      13'b1011010101000:
        _o_sv = 15'b111001011000101;
      13'b1011010101001:
        _o_sv = 15'b111001011001000;
      13'b1011010101010:
        _o_sv = 15'b111001011001010;
      13'b1011010101011:
        _o_sv = 15'b111001011001101;
      13'b1011010101100:
        _o_sv = 15'b111001011010000;
      13'b1011010101101:
        _o_sv = 15'b111001011010011;
      13'b1011010101110:
        _o_sv = 15'b111001011010101;
      13'b1011010101111:
        _o_sv = 15'b111001011011000;
      13'b1011010110000:
        _o_sv = 15'b111001011011011;
      13'b1011010110001:
        _o_sv = 15'b111001011011110;
      13'b1011010110010:
        _o_sv = 15'b111001011100001;
      13'b1011010110011:
        _o_sv = 15'b111001011100011;
      13'b1011010110100:
        _o_sv = 15'b111001011100110;
      13'b1011010110101:
        _o_sv = 15'b111001011101001;
      13'b1011010110110:
        _o_sv = 15'b111001011101100;
      13'b1011010110111:
        _o_sv = 15'b111001011101110;
      13'b1011010111000:
        _o_sv = 15'b111001011110001;
      13'b1011010111001:
        _o_sv = 15'b111001011110100;
      13'b1011010111010:
        _o_sv = 15'b111001011110111;
      13'b1011010111011:
        _o_sv = 15'b111001011111001;
      13'b1011010111100:
        _o_sv = 15'b111001011111100;
      13'b1011010111101:
        _o_sv = 15'b111001011111111;
      13'b1011010111110:
        _o_sv = 15'b111001100000010;
      13'b1011010111111:
        _o_sv = 15'b111001100000101;
      13'b1011011000000:
        _o_sv = 15'b111001100000111;
      13'b1011011000001:
        _o_sv = 15'b111001100001010;
      13'b1011011000010:
        _o_sv = 15'b111001100001101;
      13'b1011011000011:
        _o_sv = 15'b111001100010000;
      13'b1011011000100:
        _o_sv = 15'b111001100010010;
      13'b1011011000101:
        _o_sv = 15'b111001100010101;
      13'b1011011000110:
        _o_sv = 15'b111001100011000;
      13'b1011011000111:
        _o_sv = 15'b111001100011011;
      13'b1011011001000:
        _o_sv = 15'b111001100011101;
      13'b1011011001001:
        _o_sv = 15'b111001100100000;
      13'b1011011001010:
        _o_sv = 15'b111001100100011;
      13'b1011011001011:
        _o_sv = 15'b111001100100110;
      13'b1011011001100:
        _o_sv = 15'b111001100101000;
      13'b1011011001101:
        _o_sv = 15'b111001100101011;
      13'b1011011001110:
        _o_sv = 15'b111001100101110;
      13'b1011011001111:
        _o_sv = 15'b111001100110000;
      13'b1011011010000:
        _o_sv = 15'b111001100110011;
      13'b1011011010001:
        _o_sv = 15'b111001100110110;
      13'b1011011010010:
        _o_sv = 15'b111001100111001;
      13'b1011011010011:
        _o_sv = 15'b111001100111011;
      13'b1011011010100:
        _o_sv = 15'b111001100111110;
      13'b1011011010101:
        _o_sv = 15'b111001101000001;
      13'b1011011010110:
        _o_sv = 15'b111001101000100;
      13'b1011011010111:
        _o_sv = 15'b111001101000110;
      13'b1011011011000:
        _o_sv = 15'b111001101001001;
      13'b1011011011001:
        _o_sv = 15'b111001101001100;
      13'b1011011011010:
        _o_sv = 15'b111001101001111;
      13'b1011011011011:
        _o_sv = 15'b111001101010001;
      13'b1011011011100:
        _o_sv = 15'b111001101010100;
      13'b1011011011101:
        _o_sv = 15'b111001101010111;
      13'b1011011011110:
        _o_sv = 15'b111001101011001;
      13'b1011011011111:
        _o_sv = 15'b111001101011100;
      13'b1011011100000:
        _o_sv = 15'b111001101011111;
      13'b1011011100001:
        _o_sv = 15'b111001101100010;
      13'b1011011100010:
        _o_sv = 15'b111001101100100;
      13'b1011011100011:
        _o_sv = 15'b111001101100111;
      13'b1011011100100:
        _o_sv = 15'b111001101101010;
      13'b1011011100101:
        _o_sv = 15'b111001101101100;
      13'b1011011100110:
        _o_sv = 15'b111001101101111;
      13'b1011011100111:
        _o_sv = 15'b111001101110010;
      13'b1011011101000:
        _o_sv = 15'b111001101110101;
      13'b1011011101001:
        _o_sv = 15'b111001101110111;
      13'b1011011101010:
        _o_sv = 15'b111001101111010;
      13'b1011011101011:
        _o_sv = 15'b111001101111101;
      13'b1011011101100:
        _o_sv = 15'b111001101111111;
      13'b1011011101101:
        _o_sv = 15'b111001110000010;
      13'b1011011101110:
        _o_sv = 15'b111001110000101;
      13'b1011011101111:
        _o_sv = 15'b111001110001000;
      13'b1011011110000:
        _o_sv = 15'b111001110001010;
      13'b1011011110001:
        _o_sv = 15'b111001110001101;
      13'b1011011110010:
        _o_sv = 15'b111001110010000;
      13'b1011011110011:
        _o_sv = 15'b111001110010010;
      13'b1011011110100:
        _o_sv = 15'b111001110010101;
      13'b1011011110101:
        _o_sv = 15'b111001110011000;
      13'b1011011110110:
        _o_sv = 15'b111001110011011;
      13'b1011011110111:
        _o_sv = 15'b111001110011101;
      13'b1011011111000:
        _o_sv = 15'b111001110100000;
      13'b1011011111001:
        _o_sv = 15'b111001110100011;
      13'b1011011111010:
        _o_sv = 15'b111001110100101;
      13'b1011011111011:
        _o_sv = 15'b111001110101000;
      13'b1011011111100:
        _o_sv = 15'b111001110101011;
      13'b1011011111101:
        _o_sv = 15'b111001110101101;
      13'b1011011111110:
        _o_sv = 15'b111001110110000;
      13'b1011011111111:
        _o_sv = 15'b111001110110011;
      13'b1011100000000:
        _o_sv = 15'b111001110110101;
      13'b1011100000001:
        _o_sv = 15'b111001110111000;
      13'b1011100000010:
        _o_sv = 15'b111001110111011;
      13'b1011100000011:
        _o_sv = 15'b111001110111101;
      13'b1011100000100:
        _o_sv = 15'b111001111000000;
      13'b1011100000101:
        _o_sv = 15'b111001111000011;
      13'b1011100000110:
        _o_sv = 15'b111001111000110;
      13'b1011100000111:
        _o_sv = 15'b111001111001000;
      13'b1011100001000:
        _o_sv = 15'b111001111001011;
      13'b1011100001001:
        _o_sv = 15'b111001111001110;
      13'b1011100001010:
        _o_sv = 15'b111001111010000;
      13'b1011100001011:
        _o_sv = 15'b111001111010011;
      13'b1011100001100:
        _o_sv = 15'b111001111010110;
      13'b1011100001101:
        _o_sv = 15'b111001111011000;
      13'b1011100001110:
        _o_sv = 15'b111001111011011;
      13'b1011100001111:
        _o_sv = 15'b111001111011110;
      13'b1011100010000:
        _o_sv = 15'b111001111100000;
      13'b1011100010001:
        _o_sv = 15'b111001111100011;
      13'b1011100010010:
        _o_sv = 15'b111001111100110;
      13'b1011100010011:
        _o_sv = 15'b111001111101000;
      13'b1011100010100:
        _o_sv = 15'b111001111101011;
      13'b1011100010101:
        _o_sv = 15'b111001111101110;
      13'b1011100010110:
        _o_sv = 15'b111001111110000;
      13'b1011100010111:
        _o_sv = 15'b111001111110011;
      13'b1011100011000:
        _o_sv = 15'b111001111110110;
      13'b1011100011001:
        _o_sv = 15'b111001111111000;
      13'b1011100011010:
        _o_sv = 15'b111001111111011;
      13'b1011100011011:
        _o_sv = 15'b111001111111110;
      13'b1011100011100:
        _o_sv = 15'b111010000000000;
      13'b1011100011101:
        _o_sv = 15'b111010000000011;
      13'b1011100011110:
        _o_sv = 15'b111010000000110;
      13'b1011100011111:
        _o_sv = 15'b111010000001000;
      13'b1011100100000:
        _o_sv = 15'b111010000001011;
      13'b1011100100001:
        _o_sv = 15'b111010000001101;
      13'b1011100100010:
        _o_sv = 15'b111010000010000;
      13'b1011100100011:
        _o_sv = 15'b111010000010011;
      13'b1011100100100:
        _o_sv = 15'b111010000010101;
      13'b1011100100101:
        _o_sv = 15'b111010000011000;
      13'b1011100100110:
        _o_sv = 15'b111010000011011;
      13'b1011100100111:
        _o_sv = 15'b111010000011101;
      13'b1011100101000:
        _o_sv = 15'b111010000100000;
      13'b1011100101001:
        _o_sv = 15'b111010000100011;
      13'b1011100101010:
        _o_sv = 15'b111010000100101;
      13'b1011100101011:
        _o_sv = 15'b111010000101000;
      13'b1011100101100:
        _o_sv = 15'b111010000101011;
      13'b1011100101101:
        _o_sv = 15'b111010000101101;
      13'b1011100101110:
        _o_sv = 15'b111010000110000;
      13'b1011100101111:
        _o_sv = 15'b111010000110010;
      13'b1011100110000:
        _o_sv = 15'b111010000110101;
      13'b1011100110001:
        _o_sv = 15'b111010000111000;
      13'b1011100110010:
        _o_sv = 15'b111010000111010;
      13'b1011100110011:
        _o_sv = 15'b111010000111101;
      13'b1011100110100:
        _o_sv = 15'b111010001000000;
      13'b1011100110101:
        _o_sv = 15'b111010001000010;
      13'b1011100110110:
        _o_sv = 15'b111010001000101;
      13'b1011100110111:
        _o_sv = 15'b111010001001000;
      13'b1011100111000:
        _o_sv = 15'b111010001001010;
      13'b1011100111001:
        _o_sv = 15'b111010001001101;
      13'b1011100111010:
        _o_sv = 15'b111010001001111;
      13'b1011100111011:
        _o_sv = 15'b111010001010010;
      13'b1011100111100:
        _o_sv = 15'b111010001010101;
      13'b1011100111101:
        _o_sv = 15'b111010001010111;
      13'b1011100111110:
        _o_sv = 15'b111010001011010;
      13'b1011100111111:
        _o_sv = 15'b111010001011100;
      13'b1011101000000:
        _o_sv = 15'b111010001011111;
      13'b1011101000001:
        _o_sv = 15'b111010001100010;
      13'b1011101000010:
        _o_sv = 15'b111010001100100;
      13'b1011101000011:
        _o_sv = 15'b111010001100111;
      13'b1011101000100:
        _o_sv = 15'b111010001101010;
      13'b1011101000101:
        _o_sv = 15'b111010001101100;
      13'b1011101000110:
        _o_sv = 15'b111010001101111;
      13'b1011101000111:
        _o_sv = 15'b111010001110001;
      13'b1011101001000:
        _o_sv = 15'b111010001110100;
      13'b1011101001001:
        _o_sv = 15'b111010001110111;
      13'b1011101001010:
        _o_sv = 15'b111010001111001;
      13'b1011101001011:
        _o_sv = 15'b111010001111100;
      13'b1011101001100:
        _o_sv = 15'b111010001111110;
      13'b1011101001101:
        _o_sv = 15'b111010010000001;
      13'b1011101001110:
        _o_sv = 15'b111010010000100;
      13'b1011101001111:
        _o_sv = 15'b111010010000110;
      13'b1011101010000:
        _o_sv = 15'b111010010001001;
      13'b1011101010001:
        _o_sv = 15'b111010010001011;
      13'b1011101010010:
        _o_sv = 15'b111010010001110;
      13'b1011101010011:
        _o_sv = 15'b111010010010001;
      13'b1011101010100:
        _o_sv = 15'b111010010010011;
      13'b1011101010101:
        _o_sv = 15'b111010010010110;
      13'b1011101010110:
        _o_sv = 15'b111010010011000;
      13'b1011101010111:
        _o_sv = 15'b111010010011011;
      13'b1011101011000:
        _o_sv = 15'b111010010011110;
      13'b1011101011001:
        _o_sv = 15'b111010010100000;
      13'b1011101011010:
        _o_sv = 15'b111010010100011;
      13'b1011101011011:
        _o_sv = 15'b111010010100101;
      13'b1011101011100:
        _o_sv = 15'b111010010101000;
      13'b1011101011101:
        _o_sv = 15'b111010010101011;
      13'b1011101011110:
        _o_sv = 15'b111010010101101;
      13'b1011101011111:
        _o_sv = 15'b111010010110000;
      13'b1011101100000:
        _o_sv = 15'b111010010110010;
      13'b1011101100001:
        _o_sv = 15'b111010010110101;
      13'b1011101100010:
        _o_sv = 15'b111010010110111;
      13'b1011101100011:
        _o_sv = 15'b111010010111010;
      13'b1011101100100:
        _o_sv = 15'b111010010111101;
      13'b1011101100101:
        _o_sv = 15'b111010010111111;
      13'b1011101100110:
        _o_sv = 15'b111010011000010;
      13'b1011101100111:
        _o_sv = 15'b111010011000100;
      13'b1011101101000:
        _o_sv = 15'b111010011000111;
      13'b1011101101001:
        _o_sv = 15'b111010011001001;
      13'b1011101101010:
        _o_sv = 15'b111010011001100;
      13'b1011101101011:
        _o_sv = 15'b111010011001111;
      13'b1011101101100:
        _o_sv = 15'b111010011010001;
      13'b1011101101101:
        _o_sv = 15'b111010011010100;
      13'b1011101101110:
        _o_sv = 15'b111010011010110;
      13'b1011101101111:
        _o_sv = 15'b111010011011001;
      13'b1011101110000:
        _o_sv = 15'b111010011011011;
      13'b1011101110001:
        _o_sv = 15'b111010011011110;
      13'b1011101110010:
        _o_sv = 15'b111010011100001;
      13'b1011101110011:
        _o_sv = 15'b111010011100011;
      13'b1011101110100:
        _o_sv = 15'b111010011100110;
      13'b1011101110101:
        _o_sv = 15'b111010011101000;
      13'b1011101110110:
        _o_sv = 15'b111010011101011;
      13'b1011101110111:
        _o_sv = 15'b111010011101101;
      13'b1011101111000:
        _o_sv = 15'b111010011110000;
      13'b1011101111001:
        _o_sv = 15'b111010011110010;
      13'b1011101111010:
        _o_sv = 15'b111010011110101;
      13'b1011101111011:
        _o_sv = 15'b111010011111000;
      13'b1011101111100:
        _o_sv = 15'b111010011111010;
      13'b1011101111101:
        _o_sv = 15'b111010011111101;
      13'b1011101111110:
        _o_sv = 15'b111010011111111;
      13'b1011101111111:
        _o_sv = 15'b111010100000010;
      13'b1011110000000:
        _o_sv = 15'b111010100000100;
      13'b1011110000001:
        _o_sv = 15'b111010100000111;
      13'b1011110000010:
        _o_sv = 15'b111010100001001;
      13'b1011110000011:
        _o_sv = 15'b111010100001100;
      13'b1011110000100:
        _o_sv = 15'b111010100001111;
      13'b1011110000101:
        _o_sv = 15'b111010100010001;
      13'b1011110000110:
        _o_sv = 15'b111010100010100;
      13'b1011110000111:
        _o_sv = 15'b111010100010110;
      13'b1011110001000:
        _o_sv = 15'b111010100011001;
      13'b1011110001001:
        _o_sv = 15'b111010100011011;
      13'b1011110001010:
        _o_sv = 15'b111010100011110;
      13'b1011110001011:
        _o_sv = 15'b111010100100000;
      13'b1011110001100:
        _o_sv = 15'b111010100100011;
      13'b1011110001101:
        _o_sv = 15'b111010100100101;
      13'b1011110001110:
        _o_sv = 15'b111010100101000;
      13'b1011110001111:
        _o_sv = 15'b111010100101010;
      13'b1011110010000:
        _o_sv = 15'b111010100101101;
      13'b1011110010001:
        _o_sv = 15'b111010100101111;
      13'b1011110010010:
        _o_sv = 15'b111010100110010;
      13'b1011110010011:
        _o_sv = 15'b111010100110101;
      13'b1011110010100:
        _o_sv = 15'b111010100110111;
      13'b1011110010101:
        _o_sv = 15'b111010100111010;
      13'b1011110010110:
        _o_sv = 15'b111010100111100;
      13'b1011110010111:
        _o_sv = 15'b111010100111111;
      13'b1011110011000:
        _o_sv = 15'b111010101000001;
      13'b1011110011001:
        _o_sv = 15'b111010101000100;
      13'b1011110011010:
        _o_sv = 15'b111010101000110;
      13'b1011110011011:
        _o_sv = 15'b111010101001001;
      13'b1011110011100:
        _o_sv = 15'b111010101001011;
      13'b1011110011101:
        _o_sv = 15'b111010101001110;
      13'b1011110011110:
        _o_sv = 15'b111010101010000;
      13'b1011110011111:
        _o_sv = 15'b111010101010011;
      13'b1011110100000:
        _o_sv = 15'b111010101010101;
      13'b1011110100001:
        _o_sv = 15'b111010101011000;
      13'b1011110100010:
        _o_sv = 15'b111010101011010;
      13'b1011110100011:
        _o_sv = 15'b111010101011101;
      13'b1011110100100:
        _o_sv = 15'b111010101011111;
      13'b1011110100101:
        _o_sv = 15'b111010101100010;
      13'b1011110100110:
        _o_sv = 15'b111010101100100;
      13'b1011110100111:
        _o_sv = 15'b111010101100111;
      13'b1011110101000:
        _o_sv = 15'b111010101101001;
      13'b1011110101001:
        _o_sv = 15'b111010101101100;
      13'b1011110101010:
        _o_sv = 15'b111010101101110;
      13'b1011110101011:
        _o_sv = 15'b111010101110001;
      13'b1011110101100:
        _o_sv = 15'b111010101110011;
      13'b1011110101101:
        _o_sv = 15'b111010101110110;
      13'b1011110101110:
        _o_sv = 15'b111010101111000;
      13'b1011110101111:
        _o_sv = 15'b111010101111011;
      13'b1011110110000:
        _o_sv = 15'b111010101111101;
      13'b1011110110001:
        _o_sv = 15'b111010110000000;
      13'b1011110110010:
        _o_sv = 15'b111010110000010;
      13'b1011110110011:
        _o_sv = 15'b111010110000101;
      13'b1011110110100:
        _o_sv = 15'b111010110000111;
      13'b1011110110101:
        _o_sv = 15'b111010110001010;
      13'b1011110110110:
        _o_sv = 15'b111010110001100;
      13'b1011110110111:
        _o_sv = 15'b111010110001111;
      13'b1011110111000:
        _o_sv = 15'b111010110010001;
      13'b1011110111001:
        _o_sv = 15'b111010110010100;
      13'b1011110111010:
        _o_sv = 15'b111010110010110;
      13'b1011110111011:
        _o_sv = 15'b111010110011001;
      13'b1011110111100:
        _o_sv = 15'b111010110011011;
      13'b1011110111101:
        _o_sv = 15'b111010110011110;
      13'b1011110111110:
        _o_sv = 15'b111010110100000;
      13'b1011110111111:
        _o_sv = 15'b111010110100011;
      13'b1011111000000:
        _o_sv = 15'b111010110100101;
      13'b1011111000001:
        _o_sv = 15'b111010110100111;
      13'b1011111000010:
        _o_sv = 15'b111010110101010;
      13'b1011111000011:
        _o_sv = 15'b111010110101100;
      13'b1011111000100:
        _o_sv = 15'b111010110101111;
      13'b1011111000101:
        _o_sv = 15'b111010110110001;
      13'b1011111000110:
        _o_sv = 15'b111010110110100;
      13'b1011111000111:
        _o_sv = 15'b111010110110110;
      13'b1011111001000:
        _o_sv = 15'b111010110111001;
      13'b1011111001001:
        _o_sv = 15'b111010110111011;
      13'b1011111001010:
        _o_sv = 15'b111010110111110;
      13'b1011111001011:
        _o_sv = 15'b111010111000000;
      13'b1011111001100:
        _o_sv = 15'b111010111000011;
      13'b1011111001101:
        _o_sv = 15'b111010111000101;
      13'b1011111001110:
        _o_sv = 15'b111010111001000;
      13'b1011111001111:
        _o_sv = 15'b111010111001010;
      13'b1011111010000:
        _o_sv = 15'b111010111001100;
      13'b1011111010001:
        _o_sv = 15'b111010111001111;
      13'b1011111010010:
        _o_sv = 15'b111010111010001;
      13'b1011111010011:
        _o_sv = 15'b111010111010100;
      13'b1011111010100:
        _o_sv = 15'b111010111010110;
      13'b1011111010101:
        _o_sv = 15'b111010111011001;
      13'b1011111010110:
        _o_sv = 15'b111010111011011;
      13'b1011111010111:
        _o_sv = 15'b111010111011110;
      13'b1011111011000:
        _o_sv = 15'b111010111100000;
      13'b1011111011001:
        _o_sv = 15'b111010111100011;
      13'b1011111011010:
        _o_sv = 15'b111010111100101;
      13'b1011111011011:
        _o_sv = 15'b111010111100111;
      13'b1011111011100:
        _o_sv = 15'b111010111101010;
      13'b1011111011101:
        _o_sv = 15'b111010111101100;
      13'b1011111011110:
        _o_sv = 15'b111010111101111;
      13'b1011111011111:
        _o_sv = 15'b111010111110001;
      13'b1011111100000:
        _o_sv = 15'b111010111110100;
      13'b1011111100001:
        _o_sv = 15'b111010111110110;
      13'b1011111100010:
        _o_sv = 15'b111010111111001;
      13'b1011111100011:
        _o_sv = 15'b111010111111011;
      13'b1011111100100:
        _o_sv = 15'b111010111111101;
      13'b1011111100101:
        _o_sv = 15'b111011000000000;
      13'b1011111100110:
        _o_sv = 15'b111011000000010;
      13'b1011111100111:
        _o_sv = 15'b111011000000101;
      13'b1011111101000:
        _o_sv = 15'b111011000000111;
      13'b1011111101001:
        _o_sv = 15'b111011000001010;
      13'b1011111101010:
        _o_sv = 15'b111011000001100;
      13'b1011111101011:
        _o_sv = 15'b111011000001110;
      13'b1011111101100:
        _o_sv = 15'b111011000010001;
      13'b1011111101101:
        _o_sv = 15'b111011000010011;
      13'b1011111101110:
        _o_sv = 15'b111011000010110;
      13'b1011111101111:
        _o_sv = 15'b111011000011000;
      13'b1011111110000:
        _o_sv = 15'b111011000011011;
      13'b1011111110001:
        _o_sv = 15'b111011000011101;
      13'b1011111110010:
        _o_sv = 15'b111011000011111;
      13'b1011111110011:
        _o_sv = 15'b111011000100010;
      13'b1011111110100:
        _o_sv = 15'b111011000100100;
      13'b1011111110101:
        _o_sv = 15'b111011000100111;
      13'b1011111110110:
        _o_sv = 15'b111011000101001;
      13'b1011111110111:
        _o_sv = 15'b111011000101011;
      13'b1011111111000:
        _o_sv = 15'b111011000101110;
      13'b1011111111001:
        _o_sv = 15'b111011000110000;
      13'b1011111111010:
        _o_sv = 15'b111011000110011;
      13'b1011111111011:
        _o_sv = 15'b111011000110101;
      13'b1011111111100:
        _o_sv = 15'b111011000111000;
      13'b1011111111101:
        _o_sv = 15'b111011000111010;
      13'b1011111111110:
        _o_sv = 15'b111011000111100;
      13'b1011111111111:
        _o_sv = 15'b111011000111111;
      13'b1100000000000:
        _o_sv = 15'b111011001000001;
      13'b1100000000001:
        _o_sv = 15'b111011001000100;
      13'b1100000000010:
        _o_sv = 15'b111011001000110;
      13'b1100000000011:
        _o_sv = 15'b111011001001000;
      13'b1100000000100:
        _o_sv = 15'b111011001001011;
      13'b1100000000101:
        _o_sv = 15'b111011001001101;
      13'b1100000000110:
        _o_sv = 15'b111011001010000;
      13'b1100000000111:
        _o_sv = 15'b111011001010010;
      13'b1100000001000:
        _o_sv = 15'b111011001010100;
      13'b1100000001001:
        _o_sv = 15'b111011001010111;
      13'b1100000001010:
        _o_sv = 15'b111011001011001;
      13'b1100000001011:
        _o_sv = 15'b111011001011100;
      13'b1100000001100:
        _o_sv = 15'b111011001011110;
      13'b1100000001101:
        _o_sv = 15'b111011001100000;
      13'b1100000001110:
        _o_sv = 15'b111011001100011;
      13'b1100000001111:
        _o_sv = 15'b111011001100101;
      13'b1100000010000:
        _o_sv = 15'b111011001101000;
      13'b1100000010001:
        _o_sv = 15'b111011001101010;
      13'b1100000010010:
        _o_sv = 15'b111011001101100;
      13'b1100000010011:
        _o_sv = 15'b111011001101111;
      13'b1100000010100:
        _o_sv = 15'b111011001110001;
      13'b1100000010101:
        _o_sv = 15'b111011001110011;
      13'b1100000010110:
        _o_sv = 15'b111011001110110;
      13'b1100000010111:
        _o_sv = 15'b111011001111000;
      13'b1100000011000:
        _o_sv = 15'b111011001111011;
      13'b1100000011001:
        _o_sv = 15'b111011001111101;
      13'b1100000011010:
        _o_sv = 15'b111011001111111;
      13'b1100000011011:
        _o_sv = 15'b111011010000010;
      13'b1100000011100:
        _o_sv = 15'b111011010000100;
      13'b1100000011101:
        _o_sv = 15'b111011010000110;
      13'b1100000011110:
        _o_sv = 15'b111011010001001;
      13'b1100000011111:
        _o_sv = 15'b111011010001011;
      13'b1100000100000:
        _o_sv = 15'b111011010001110;
      13'b1100000100001:
        _o_sv = 15'b111011010010000;
      13'b1100000100010:
        _o_sv = 15'b111011010010010;
      13'b1100000100011:
        _o_sv = 15'b111011010010101;
      13'b1100000100100:
        _o_sv = 15'b111011010010111;
      13'b1100000100101:
        _o_sv = 15'b111011010011001;
      13'b1100000100110:
        _o_sv = 15'b111011010011100;
      13'b1100000100111:
        _o_sv = 15'b111011010011110;
      13'b1100000101000:
        _o_sv = 15'b111011010100000;
      13'b1100000101001:
        _o_sv = 15'b111011010100011;
      13'b1100000101010:
        _o_sv = 15'b111011010100101;
      13'b1100000101011:
        _o_sv = 15'b111011010101000;
      13'b1100000101100:
        _o_sv = 15'b111011010101010;
      13'b1100000101101:
        _o_sv = 15'b111011010101100;
      13'b1100000101110:
        _o_sv = 15'b111011010101111;
      13'b1100000101111:
        _o_sv = 15'b111011010110001;
      13'b1100000110000:
        _o_sv = 15'b111011010110011;
      13'b1100000110001:
        _o_sv = 15'b111011010110110;
      13'b1100000110010:
        _o_sv = 15'b111011010111000;
      13'b1100000110011:
        _o_sv = 15'b111011010111010;
      13'b1100000110100:
        _o_sv = 15'b111011010111101;
      13'b1100000110101:
        _o_sv = 15'b111011010111111;
      13'b1100000110110:
        _o_sv = 15'b111011011000001;
      13'b1100000110111:
        _o_sv = 15'b111011011000100;
      13'b1100000111000:
        _o_sv = 15'b111011011000110;
      13'b1100000111001:
        _o_sv = 15'b111011011001000;
      13'b1100000111010:
        _o_sv = 15'b111011011001011;
      13'b1100000111011:
        _o_sv = 15'b111011011001101;
      13'b1100000111100:
        _o_sv = 15'b111011011001111;
      13'b1100000111101:
        _o_sv = 15'b111011011010010;
      13'b1100000111110:
        _o_sv = 15'b111011011010100;
      13'b1100000111111:
        _o_sv = 15'b111011011010110;
      13'b1100001000000:
        _o_sv = 15'b111011011011001;
      13'b1100001000001:
        _o_sv = 15'b111011011011011;
      13'b1100001000010:
        _o_sv = 15'b111011011011101;
      13'b1100001000011:
        _o_sv = 15'b111011011100000;
      13'b1100001000100:
        _o_sv = 15'b111011011100010;
      13'b1100001000101:
        _o_sv = 15'b111011011100100;
      13'b1100001000110:
        _o_sv = 15'b111011011100111;
      13'b1100001000111:
        _o_sv = 15'b111011011101001;
      13'b1100001001000:
        _o_sv = 15'b111011011101011;
      13'b1100001001001:
        _o_sv = 15'b111011011101110;
      13'b1100001001010:
        _o_sv = 15'b111011011110000;
      13'b1100001001011:
        _o_sv = 15'b111011011110010;
      13'b1100001001100:
        _o_sv = 15'b111011011110101;
      13'b1100001001101:
        _o_sv = 15'b111011011110111;
      13'b1100001001110:
        _o_sv = 15'b111011011111001;
      13'b1100001001111:
        _o_sv = 15'b111011011111100;
      13'b1100001010000:
        _o_sv = 15'b111011011111110;
      13'b1100001010001:
        _o_sv = 15'b111011100000000;
      13'b1100001010010:
        _o_sv = 15'b111011100000011;
      13'b1100001010011:
        _o_sv = 15'b111011100000101;
      13'b1100001010100:
        _o_sv = 15'b111011100000111;
      13'b1100001010101:
        _o_sv = 15'b111011100001010;
      13'b1100001010110:
        _o_sv = 15'b111011100001100;
      13'b1100001010111:
        _o_sv = 15'b111011100001110;
      13'b1100001011000:
        _o_sv = 15'b111011100010000;
      13'b1100001011001:
        _o_sv = 15'b111011100010011;
      13'b1100001011010:
        _o_sv = 15'b111011100010101;
      13'b1100001011011:
        _o_sv = 15'b111011100010111;
      13'b1100001011100:
        _o_sv = 15'b111011100011010;
      13'b1100001011101:
        _o_sv = 15'b111011100011100;
      13'b1100001011110:
        _o_sv = 15'b111011100011110;
      13'b1100001011111:
        _o_sv = 15'b111011100100001;
      13'b1100001100000:
        _o_sv = 15'b111011100100011;
      13'b1100001100001:
        _o_sv = 15'b111011100100101;
      13'b1100001100010:
        _o_sv = 15'b111011100100111;
      13'b1100001100011:
        _o_sv = 15'b111011100101010;
      13'b1100001100100:
        _o_sv = 15'b111011100101100;
      13'b1100001100101:
        _o_sv = 15'b111011100101110;
      13'b1100001100110:
        _o_sv = 15'b111011100110001;
      13'b1100001100111:
        _o_sv = 15'b111011100110011;
      13'b1100001101000:
        _o_sv = 15'b111011100110101;
      13'b1100001101001:
        _o_sv = 15'b111011100111000;
      13'b1100001101010:
        _o_sv = 15'b111011100111010;
      13'b1100001101011:
        _o_sv = 15'b111011100111100;
      13'b1100001101100:
        _o_sv = 15'b111011100111110;
      13'b1100001101101:
        _o_sv = 15'b111011101000001;
      13'b1100001101110:
        _o_sv = 15'b111011101000011;
      13'b1100001101111:
        _o_sv = 15'b111011101000101;
      13'b1100001110000:
        _o_sv = 15'b111011101000111;
      13'b1100001110001:
        _o_sv = 15'b111011101001010;
      13'b1100001110010:
        _o_sv = 15'b111011101001100;
      13'b1100001110011:
        _o_sv = 15'b111011101001110;
      13'b1100001110100:
        _o_sv = 15'b111011101010001;
      13'b1100001110101:
        _o_sv = 15'b111011101010011;
      13'b1100001110110:
        _o_sv = 15'b111011101010101;
      13'b1100001110111:
        _o_sv = 15'b111011101010111;
      13'b1100001111000:
        _o_sv = 15'b111011101011010;
      13'b1100001111001:
        _o_sv = 15'b111011101011100;
      13'b1100001111010:
        _o_sv = 15'b111011101011110;
      13'b1100001111011:
        _o_sv = 15'b111011101100000;
      13'b1100001111100:
        _o_sv = 15'b111011101100011;
      13'b1100001111101:
        _o_sv = 15'b111011101100101;
      13'b1100001111110:
        _o_sv = 15'b111011101100111;
      13'b1100001111111:
        _o_sv = 15'b111011101101010;
      13'b1100010000000:
        _o_sv = 15'b111011101101100;
      13'b1100010000001:
        _o_sv = 15'b111011101101110;
      13'b1100010000010:
        _o_sv = 15'b111011101110000;
      13'b1100010000011:
        _o_sv = 15'b111011101110011;
      13'b1100010000100:
        _o_sv = 15'b111011101110101;
      13'b1100010000101:
        _o_sv = 15'b111011101110111;
      13'b1100010000110:
        _o_sv = 15'b111011101111001;
      13'b1100010000111:
        _o_sv = 15'b111011101111100;
      13'b1100010001000:
        _o_sv = 15'b111011101111110;
      13'b1100010001001:
        _o_sv = 15'b111011110000000;
      13'b1100010001010:
        _o_sv = 15'b111011110000010;
      13'b1100010001011:
        _o_sv = 15'b111011110000101;
      13'b1100010001100:
        _o_sv = 15'b111011110000111;
      13'b1100010001101:
        _o_sv = 15'b111011110001001;
      13'b1100010001110:
        _o_sv = 15'b111011110001011;
      13'b1100010001111:
        _o_sv = 15'b111011110001110;
      13'b1100010010000:
        _o_sv = 15'b111011110010000;
      13'b1100010010001:
        _o_sv = 15'b111011110010010;
      13'b1100010010010:
        _o_sv = 15'b111011110010100;
      13'b1100010010011:
        _o_sv = 15'b111011110010111;
      13'b1100010010100:
        _o_sv = 15'b111011110011001;
      13'b1100010010101:
        _o_sv = 15'b111011110011011;
      13'b1100010010110:
        _o_sv = 15'b111011110011101;
      13'b1100010010111:
        _o_sv = 15'b111011110100000;
      13'b1100010011000:
        _o_sv = 15'b111011110100010;
      13'b1100010011001:
        _o_sv = 15'b111011110100100;
      13'b1100010011010:
        _o_sv = 15'b111011110100110;
      13'b1100010011011:
        _o_sv = 15'b111011110101000;
      13'b1100010011100:
        _o_sv = 15'b111011110101011;
      13'b1100010011101:
        _o_sv = 15'b111011110101101;
      13'b1100010011110:
        _o_sv = 15'b111011110101111;
      13'b1100010011111:
        _o_sv = 15'b111011110110001;
      13'b1100010100000:
        _o_sv = 15'b111011110110100;
      13'b1100010100001:
        _o_sv = 15'b111011110110110;
      13'b1100010100010:
        _o_sv = 15'b111011110111000;
      13'b1100010100011:
        _o_sv = 15'b111011110111010;
      13'b1100010100100:
        _o_sv = 15'b111011110111100;
      13'b1100010100101:
        _o_sv = 15'b111011110111111;
      13'b1100010100110:
        _o_sv = 15'b111011111000001;
      13'b1100010100111:
        _o_sv = 15'b111011111000011;
      13'b1100010101000:
        _o_sv = 15'b111011111000101;
      13'b1100010101001:
        _o_sv = 15'b111011111001000;
      13'b1100010101010:
        _o_sv = 15'b111011111001010;
      13'b1100010101011:
        _o_sv = 15'b111011111001100;
      13'b1100010101100:
        _o_sv = 15'b111011111001110;
      13'b1100010101101:
        _o_sv = 15'b111011111010000;
      13'b1100010101110:
        _o_sv = 15'b111011111010011;
      13'b1100010101111:
        _o_sv = 15'b111011111010101;
      13'b1100010110000:
        _o_sv = 15'b111011111010111;
      13'b1100010110001:
        _o_sv = 15'b111011111011001;
      13'b1100010110010:
        _o_sv = 15'b111011111011011;
      13'b1100010110011:
        _o_sv = 15'b111011111011110;
      13'b1100010110100:
        _o_sv = 15'b111011111100000;
      13'b1100010110101:
        _o_sv = 15'b111011111100010;
      13'b1100010110110:
        _o_sv = 15'b111011111100100;
      13'b1100010110111:
        _o_sv = 15'b111011111100110;
      13'b1100010111000:
        _o_sv = 15'b111011111101001;
      13'b1100010111001:
        _o_sv = 15'b111011111101011;
      13'b1100010111010:
        _o_sv = 15'b111011111101101;
      13'b1100010111011:
        _o_sv = 15'b111011111101111;
      13'b1100010111100:
        _o_sv = 15'b111011111110001;
      13'b1100010111101:
        _o_sv = 15'b111011111110100;
      13'b1100010111110:
        _o_sv = 15'b111011111110110;
      13'b1100010111111:
        _o_sv = 15'b111011111111000;
      13'b1100011000000:
        _o_sv = 15'b111011111111010;
      13'b1100011000001:
        _o_sv = 15'b111011111111100;
      13'b1100011000010:
        _o_sv = 15'b111011111111111;
      13'b1100011000011:
        _o_sv = 15'b111100000000001;
      13'b1100011000100:
        _o_sv = 15'b111100000000011;
      13'b1100011000101:
        _o_sv = 15'b111100000000101;
      13'b1100011000110:
        _o_sv = 15'b111100000000111;
      13'b1100011000111:
        _o_sv = 15'b111100000001010;
      13'b1100011001000:
        _o_sv = 15'b111100000001100;
      13'b1100011001001:
        _o_sv = 15'b111100000001110;
      13'b1100011001010:
        _o_sv = 15'b111100000010000;
      13'b1100011001011:
        _o_sv = 15'b111100000010010;
      13'b1100011001100:
        _o_sv = 15'b111100000010100;
      13'b1100011001101:
        _o_sv = 15'b111100000010111;
      13'b1100011001110:
        _o_sv = 15'b111100000011001;
      13'b1100011001111:
        _o_sv = 15'b111100000011011;
      13'b1100011010000:
        _o_sv = 15'b111100000011101;
      13'b1100011010001:
        _o_sv = 15'b111100000011111;
      13'b1100011010010:
        _o_sv = 15'b111100000100001;
      13'b1100011010011:
        _o_sv = 15'b111100000100100;
      13'b1100011010100:
        _o_sv = 15'b111100000100110;
      13'b1100011010101:
        _o_sv = 15'b111100000101000;
      13'b1100011010110:
        _o_sv = 15'b111100000101010;
      13'b1100011010111:
        _o_sv = 15'b111100000101100;
      13'b1100011011000:
        _o_sv = 15'b111100000101110;
      13'b1100011011001:
        _o_sv = 15'b111100000110001;
      13'b1100011011010:
        _o_sv = 15'b111100000110011;
      13'b1100011011011:
        _o_sv = 15'b111100000110101;
      13'b1100011011100:
        _o_sv = 15'b111100000110111;
      13'b1100011011101:
        _o_sv = 15'b111100000111001;
      13'b1100011011110:
        _o_sv = 15'b111100000111011;
      13'b1100011011111:
        _o_sv = 15'b111100000111110;
      13'b1100011100000:
        _o_sv = 15'b111100001000000;
      13'b1100011100001:
        _o_sv = 15'b111100001000010;
      13'b1100011100010:
        _o_sv = 15'b111100001000100;
      13'b1100011100011:
        _o_sv = 15'b111100001000110;
      13'b1100011100100:
        _o_sv = 15'b111100001001000;
      13'b1100011100101:
        _o_sv = 15'b111100001001010;
      13'b1100011100110:
        _o_sv = 15'b111100001001101;
      13'b1100011100111:
        _o_sv = 15'b111100001001111;
      13'b1100011101000:
        _o_sv = 15'b111100001010001;
      13'b1100011101001:
        _o_sv = 15'b111100001010011;
      13'b1100011101010:
        _o_sv = 15'b111100001010101;
      13'b1100011101011:
        _o_sv = 15'b111100001010111;
      13'b1100011101100:
        _o_sv = 15'b111100001011001;
      13'b1100011101101:
        _o_sv = 15'b111100001011100;
      13'b1100011101110:
        _o_sv = 15'b111100001011110;
      13'b1100011101111:
        _o_sv = 15'b111100001100000;
      13'b1100011110000:
        _o_sv = 15'b111100001100010;
      13'b1100011110001:
        _o_sv = 15'b111100001100100;
      13'b1100011110010:
        _o_sv = 15'b111100001100110;
      13'b1100011110011:
        _o_sv = 15'b111100001101000;
      13'b1100011110100:
        _o_sv = 15'b111100001101011;
      13'b1100011110101:
        _o_sv = 15'b111100001101101;
      13'b1100011110110:
        _o_sv = 15'b111100001101111;
      13'b1100011110111:
        _o_sv = 15'b111100001110001;
      13'b1100011111000:
        _o_sv = 15'b111100001110011;
      13'b1100011111001:
        _o_sv = 15'b111100001110101;
      13'b1100011111010:
        _o_sv = 15'b111100001110111;
      13'b1100011111011:
        _o_sv = 15'b111100001111001;
      13'b1100011111100:
        _o_sv = 15'b111100001111100;
      13'b1100011111101:
        _o_sv = 15'b111100001111110;
      13'b1100011111110:
        _o_sv = 15'b111100010000000;
      13'b1100011111111:
        _o_sv = 15'b111100010000010;
      13'b1100100000000:
        _o_sv = 15'b111100010000100;
      13'b1100100000001:
        _o_sv = 15'b111100010000110;
      13'b1100100000010:
        _o_sv = 15'b111100010001000;
      13'b1100100000011:
        _o_sv = 15'b111100010001010;
      13'b1100100000100:
        _o_sv = 15'b111100010001100;
      13'b1100100000101:
        _o_sv = 15'b111100010001111;
      13'b1100100000110:
        _o_sv = 15'b111100010010001;
      13'b1100100000111:
        _o_sv = 15'b111100010010011;
      13'b1100100001000:
        _o_sv = 15'b111100010010101;
      13'b1100100001001:
        _o_sv = 15'b111100010010111;
      13'b1100100001010:
        _o_sv = 15'b111100010011001;
      13'b1100100001011:
        _o_sv = 15'b111100010011011;
      13'b1100100001100:
        _o_sv = 15'b111100010011101;
      13'b1100100001101:
        _o_sv = 15'b111100010011111;
      13'b1100100001110:
        _o_sv = 15'b111100010100010;
      13'b1100100001111:
        _o_sv = 15'b111100010100100;
      13'b1100100010000:
        _o_sv = 15'b111100010100110;
      13'b1100100010001:
        _o_sv = 15'b111100010101000;
      13'b1100100010010:
        _o_sv = 15'b111100010101010;
      13'b1100100010011:
        _o_sv = 15'b111100010101100;
      13'b1100100010100:
        _o_sv = 15'b111100010101110;
      13'b1100100010101:
        _o_sv = 15'b111100010110000;
      13'b1100100010110:
        _o_sv = 15'b111100010110010;
      13'b1100100010111:
        _o_sv = 15'b111100010110100;
      13'b1100100011000:
        _o_sv = 15'b111100010110110;
      13'b1100100011001:
        _o_sv = 15'b111100010111001;
      13'b1100100011010:
        _o_sv = 15'b111100010111011;
      13'b1100100011011:
        _o_sv = 15'b111100010111101;
      13'b1100100011100:
        _o_sv = 15'b111100010111111;
      13'b1100100011101:
        _o_sv = 15'b111100011000001;
      13'b1100100011110:
        _o_sv = 15'b111100011000011;
      13'b1100100011111:
        _o_sv = 15'b111100011000101;
      13'b1100100100000:
        _o_sv = 15'b111100011000111;
      13'b1100100100001:
        _o_sv = 15'b111100011001001;
      13'b1100100100010:
        _o_sv = 15'b111100011001011;
      13'b1100100100011:
        _o_sv = 15'b111100011001101;
      13'b1100100100100:
        _o_sv = 15'b111100011001111;
      13'b1100100100101:
        _o_sv = 15'b111100011010010;
      13'b1100100100110:
        _o_sv = 15'b111100011010100;
      13'b1100100100111:
        _o_sv = 15'b111100011010110;
      13'b1100100101000:
        _o_sv = 15'b111100011011000;
      13'b1100100101001:
        _o_sv = 15'b111100011011010;
      13'b1100100101010:
        _o_sv = 15'b111100011011100;
      13'b1100100101011:
        _o_sv = 15'b111100011011110;
      13'b1100100101100:
        _o_sv = 15'b111100011100000;
      13'b1100100101101:
        _o_sv = 15'b111100011100010;
      13'b1100100101110:
        _o_sv = 15'b111100011100100;
      13'b1100100101111:
        _o_sv = 15'b111100011100110;
      13'b1100100110000:
        _o_sv = 15'b111100011101000;
      13'b1100100110001:
        _o_sv = 15'b111100011101010;
      13'b1100100110010:
        _o_sv = 15'b111100011101100;
      13'b1100100110011:
        _o_sv = 15'b111100011101110;
      13'b1100100110100:
        _o_sv = 15'b111100011110001;
      13'b1100100110101:
        _o_sv = 15'b111100011110011;
      13'b1100100110110:
        _o_sv = 15'b111100011110101;
      13'b1100100110111:
        _o_sv = 15'b111100011110111;
      13'b1100100111000:
        _o_sv = 15'b111100011111001;
      13'b1100100111001:
        _o_sv = 15'b111100011111011;
      13'b1100100111010:
        _o_sv = 15'b111100011111101;
      13'b1100100111011:
        _o_sv = 15'b111100011111111;
      13'b1100100111100:
        _o_sv = 15'b111100100000001;
      13'b1100100111101:
        _o_sv = 15'b111100100000011;
      13'b1100100111110:
        _o_sv = 15'b111100100000101;
      13'b1100100111111:
        _o_sv = 15'b111100100000111;
      13'b1100101000000:
        _o_sv = 15'b111100100001001;
      13'b1100101000001:
        _o_sv = 15'b111100100001011;
      13'b1100101000010:
        _o_sv = 15'b111100100001101;
      13'b1100101000011:
        _o_sv = 15'b111100100001111;
      13'b1100101000100:
        _o_sv = 15'b111100100010001;
      13'b1100101000101:
        _o_sv = 15'b111100100010011;
      13'b1100101000110:
        _o_sv = 15'b111100100010101;
      13'b1100101000111:
        _o_sv = 15'b111100100010111;
      13'b1100101001000:
        _o_sv = 15'b111100100011001;
      13'b1100101001001:
        _o_sv = 15'b111100100011100;
      13'b1100101001010:
        _o_sv = 15'b111100100011110;
      13'b1100101001011:
        _o_sv = 15'b111100100100000;
      13'b1100101001100:
        _o_sv = 15'b111100100100010;
      13'b1100101001101:
        _o_sv = 15'b111100100100100;
      13'b1100101001110:
        _o_sv = 15'b111100100100110;
      13'b1100101001111:
        _o_sv = 15'b111100100101000;
      13'b1100101010000:
        _o_sv = 15'b111100100101010;
      13'b1100101010001:
        _o_sv = 15'b111100100101100;
      13'b1100101010010:
        _o_sv = 15'b111100100101110;
      13'b1100101010011:
        _o_sv = 15'b111100100110000;
      13'b1100101010100:
        _o_sv = 15'b111100100110010;
      13'b1100101010101:
        _o_sv = 15'b111100100110100;
      13'b1100101010110:
        _o_sv = 15'b111100100110110;
      13'b1100101010111:
        _o_sv = 15'b111100100111000;
      13'b1100101011000:
        _o_sv = 15'b111100100111010;
      13'b1100101011001:
        _o_sv = 15'b111100100111100;
      13'b1100101011010:
        _o_sv = 15'b111100100111110;
      13'b1100101011011:
        _o_sv = 15'b111100101000000;
      13'b1100101011100:
        _o_sv = 15'b111100101000010;
      13'b1100101011101:
        _o_sv = 15'b111100101000100;
      13'b1100101011110:
        _o_sv = 15'b111100101000110;
      13'b1100101011111:
        _o_sv = 15'b111100101001000;
      13'b1100101100000:
        _o_sv = 15'b111100101001010;
      13'b1100101100001:
        _o_sv = 15'b111100101001100;
      13'b1100101100010:
        _o_sv = 15'b111100101001110;
      13'b1100101100011:
        _o_sv = 15'b111100101010000;
      13'b1100101100100:
        _o_sv = 15'b111100101010010;
      13'b1100101100101:
        _o_sv = 15'b111100101010100;
      13'b1100101100110:
        _o_sv = 15'b111100101010110;
      13'b1100101100111:
        _o_sv = 15'b111100101011000;
      13'b1100101101000:
        _o_sv = 15'b111100101011010;
      13'b1100101101001:
        _o_sv = 15'b111100101011100;
      13'b1100101101010:
        _o_sv = 15'b111100101011110;
      13'b1100101101011:
        _o_sv = 15'b111100101100000;
      13'b1100101101100:
        _o_sv = 15'b111100101100010;
      13'b1100101101101:
        _o_sv = 15'b111100101100100;
      13'b1100101101110:
        _o_sv = 15'b111100101100110;
      13'b1100101101111:
        _o_sv = 15'b111100101101000;
      13'b1100101110000:
        _o_sv = 15'b111100101101010;
      13'b1100101110001:
        _o_sv = 15'b111100101101100;
      13'b1100101110010:
        _o_sv = 15'b111100101101110;
      13'b1100101110011:
        _o_sv = 15'b111100101110000;
      13'b1100101110100:
        _o_sv = 15'b111100101110010;
      13'b1100101110101:
        _o_sv = 15'b111100101110100;
      13'b1100101110110:
        _o_sv = 15'b111100101110110;
      13'b1100101110111:
        _o_sv = 15'b111100101111000;
      13'b1100101111000:
        _o_sv = 15'b111100101111010;
      13'b1100101111001:
        _o_sv = 15'b111100101111100;
      13'b1100101111010:
        _o_sv = 15'b111100101111110;
      13'b1100101111011:
        _o_sv = 15'b111100110000000;
      13'b1100101111100:
        _o_sv = 15'b111100110000010;
      13'b1100101111101:
        _o_sv = 15'b111100110000100;
      13'b1100101111110:
        _o_sv = 15'b111100110000110;
      13'b1100101111111:
        _o_sv = 15'b111100110001000;
      13'b1100110000000:
        _o_sv = 15'b111100110001010;
      13'b1100110000001:
        _o_sv = 15'b111100110001100;
      13'b1100110000010:
        _o_sv = 15'b111100110001110;
      13'b1100110000011:
        _o_sv = 15'b111100110010000;
      13'b1100110000100:
        _o_sv = 15'b111100110010010;
      13'b1100110000101:
        _o_sv = 15'b111100110010011;
      13'b1100110000110:
        _o_sv = 15'b111100110010101;
      13'b1100110000111:
        _o_sv = 15'b111100110010111;
      13'b1100110001000:
        _o_sv = 15'b111100110011001;
      13'b1100110001001:
        _o_sv = 15'b111100110011011;
      13'b1100110001010:
        _o_sv = 15'b111100110011101;
      13'b1100110001011:
        _o_sv = 15'b111100110011111;
      13'b1100110001100:
        _o_sv = 15'b111100110100001;
      13'b1100110001101:
        _o_sv = 15'b111100110100011;
      13'b1100110001110:
        _o_sv = 15'b111100110100101;
      13'b1100110001111:
        _o_sv = 15'b111100110100111;
      13'b1100110010000:
        _o_sv = 15'b111100110101001;
      13'b1100110010001:
        _o_sv = 15'b111100110101011;
      13'b1100110010010:
        _o_sv = 15'b111100110101101;
      13'b1100110010011:
        _o_sv = 15'b111100110101111;
      13'b1100110010100:
        _o_sv = 15'b111100110110001;
      13'b1100110010101:
        _o_sv = 15'b111100110110011;
      13'b1100110010110:
        _o_sv = 15'b111100110110101;
      13'b1100110010111:
        _o_sv = 15'b111100110110111;
      13'b1100110011000:
        _o_sv = 15'b111100110111001;
      13'b1100110011001:
        _o_sv = 15'b111100110111011;
      13'b1100110011010:
        _o_sv = 15'b111100110111100;
      13'b1100110011011:
        _o_sv = 15'b111100110111110;
      13'b1100110011100:
        _o_sv = 15'b111100111000000;
      13'b1100110011101:
        _o_sv = 15'b111100111000010;
      13'b1100110011110:
        _o_sv = 15'b111100111000100;
      13'b1100110011111:
        _o_sv = 15'b111100111000110;
      13'b1100110100000:
        _o_sv = 15'b111100111001000;
      13'b1100110100001:
        _o_sv = 15'b111100111001010;
      13'b1100110100010:
        _o_sv = 15'b111100111001100;
      13'b1100110100011:
        _o_sv = 15'b111100111001110;
      13'b1100110100100:
        _o_sv = 15'b111100111010000;
      13'b1100110100101:
        _o_sv = 15'b111100111010010;
      13'b1100110100110:
        _o_sv = 15'b111100111010100;
      13'b1100110100111:
        _o_sv = 15'b111100111010110;
      13'b1100110101000:
        _o_sv = 15'b111100111011000;
      13'b1100110101001:
        _o_sv = 15'b111100111011001;
      13'b1100110101010:
        _o_sv = 15'b111100111011011;
      13'b1100110101011:
        _o_sv = 15'b111100111011101;
      13'b1100110101100:
        _o_sv = 15'b111100111011111;
      13'b1100110101101:
        _o_sv = 15'b111100111100001;
      13'b1100110101110:
        _o_sv = 15'b111100111100011;
      13'b1100110101111:
        _o_sv = 15'b111100111100101;
      13'b1100110110000:
        _o_sv = 15'b111100111100111;
      13'b1100110110001:
        _o_sv = 15'b111100111101001;
      13'b1100110110010:
        _o_sv = 15'b111100111101011;
      13'b1100110110011:
        _o_sv = 15'b111100111101101;
      13'b1100110110100:
        _o_sv = 15'b111100111101111;
      13'b1100110110101:
        _o_sv = 15'b111100111110000;
      13'b1100110110110:
        _o_sv = 15'b111100111110010;
      13'b1100110110111:
        _o_sv = 15'b111100111110100;
      13'b1100110111000:
        _o_sv = 15'b111100111110110;
      13'b1100110111001:
        _o_sv = 15'b111100111111000;
      13'b1100110111010:
        _o_sv = 15'b111100111111010;
      13'b1100110111011:
        _o_sv = 15'b111100111111100;
      13'b1100110111100:
        _o_sv = 15'b111100111111110;
      13'b1100110111101:
        _o_sv = 15'b111101000000000;
      13'b1100110111110:
        _o_sv = 15'b111101000000010;
      13'b1100110111111:
        _o_sv = 15'b111101000000100;
      13'b1100111000000:
        _o_sv = 15'b111101000000101;
      13'b1100111000001:
        _o_sv = 15'b111101000000111;
      13'b1100111000010:
        _o_sv = 15'b111101000001001;
      13'b1100111000011:
        _o_sv = 15'b111101000001011;
      13'b1100111000100:
        _o_sv = 15'b111101000001101;
      13'b1100111000101:
        _o_sv = 15'b111101000001111;
      13'b1100111000110:
        _o_sv = 15'b111101000010001;
      13'b1100111000111:
        _o_sv = 15'b111101000010011;
      13'b1100111001000:
        _o_sv = 15'b111101000010101;
      13'b1100111001001:
        _o_sv = 15'b111101000010110;
      13'b1100111001010:
        _o_sv = 15'b111101000011000;
      13'b1100111001011:
        _o_sv = 15'b111101000011010;
      13'b1100111001100:
        _o_sv = 15'b111101000011100;
      13'b1100111001101:
        _o_sv = 15'b111101000011110;
      13'b1100111001110:
        _o_sv = 15'b111101000100000;
      13'b1100111001111:
        _o_sv = 15'b111101000100010;
      13'b1100111010000:
        _o_sv = 15'b111101000100100;
      13'b1100111010001:
        _o_sv = 15'b111101000100110;
      13'b1100111010010:
        _o_sv = 15'b111101000100111;
      13'b1100111010011:
        _o_sv = 15'b111101000101001;
      13'b1100111010100:
        _o_sv = 15'b111101000101011;
      13'b1100111010101:
        _o_sv = 15'b111101000101101;
      13'b1100111010110:
        _o_sv = 15'b111101000101111;
      13'b1100111010111:
        _o_sv = 15'b111101000110001;
      13'b1100111011000:
        _o_sv = 15'b111101000110011;
      13'b1100111011001:
        _o_sv = 15'b111101000110101;
      13'b1100111011010:
        _o_sv = 15'b111101000110110;
      13'b1100111011011:
        _o_sv = 15'b111101000111000;
      13'b1100111011100:
        _o_sv = 15'b111101000111010;
      13'b1100111011101:
        _o_sv = 15'b111101000111100;
      13'b1100111011110:
        _o_sv = 15'b111101000111110;
      13'b1100111011111:
        _o_sv = 15'b111101001000000;
      13'b1100111100000:
        _o_sv = 15'b111101001000010;
      13'b1100111100001:
        _o_sv = 15'b111101001000011;
      13'b1100111100010:
        _o_sv = 15'b111101001000101;
      13'b1100111100011:
        _o_sv = 15'b111101001000111;
      13'b1100111100100:
        _o_sv = 15'b111101001001001;
      13'b1100111100101:
        _o_sv = 15'b111101001001011;
      13'b1100111100110:
        _o_sv = 15'b111101001001101;
      13'b1100111100111:
        _o_sv = 15'b111101001001111;
      13'b1100111101000:
        _o_sv = 15'b111101001010000;
      13'b1100111101001:
        _o_sv = 15'b111101001010010;
      13'b1100111101010:
        _o_sv = 15'b111101001010100;
      13'b1100111101011:
        _o_sv = 15'b111101001010110;
      13'b1100111101100:
        _o_sv = 15'b111101001011000;
      13'b1100111101101:
        _o_sv = 15'b111101001011010;
      13'b1100111101110:
        _o_sv = 15'b111101001011100;
      13'b1100111101111:
        _o_sv = 15'b111101001011101;
      13'b1100111110000:
        _o_sv = 15'b111101001011111;
      13'b1100111110001:
        _o_sv = 15'b111101001100001;
      13'b1100111110010:
        _o_sv = 15'b111101001100011;
      13'b1100111110011:
        _o_sv = 15'b111101001100101;
      13'b1100111110100:
        _o_sv = 15'b111101001100111;
      13'b1100111110101:
        _o_sv = 15'b111101001101000;
      13'b1100111110110:
        _o_sv = 15'b111101001101010;
      13'b1100111110111:
        _o_sv = 15'b111101001101100;
      13'b1100111111000:
        _o_sv = 15'b111101001101110;
      13'b1100111111001:
        _o_sv = 15'b111101001110000;
      13'b1100111111010:
        _o_sv = 15'b111101001110010;
      13'b1100111111011:
        _o_sv = 15'b111101001110011;
      13'b1100111111100:
        _o_sv = 15'b111101001110101;
      13'b1100111111101:
        _o_sv = 15'b111101001110111;
      13'b1100111111110:
        _o_sv = 15'b111101001111001;
      13'b1100111111111:
        _o_sv = 15'b111101001111011;
      13'b1101000000000:
        _o_sv = 15'b111101001111101;
      13'b1101000000001:
        _o_sv = 15'b111101001111110;
      13'b1101000000010:
        _o_sv = 15'b111101010000000;
      13'b1101000000011:
        _o_sv = 15'b111101010000010;
      13'b1101000000100:
        _o_sv = 15'b111101010000100;
      13'b1101000000101:
        _o_sv = 15'b111101010000110;
      13'b1101000000110:
        _o_sv = 15'b111101010000111;
      13'b1101000000111:
        _o_sv = 15'b111101010001001;
      13'b1101000001000:
        _o_sv = 15'b111101010001011;
      13'b1101000001001:
        _o_sv = 15'b111101010001101;
      13'b1101000001010:
        _o_sv = 15'b111101010001111;
      13'b1101000001011:
        _o_sv = 15'b111101010010001;
      13'b1101000001100:
        _o_sv = 15'b111101010010010;
      13'b1101000001101:
        _o_sv = 15'b111101010010100;
      13'b1101000001110:
        _o_sv = 15'b111101010010110;
      13'b1101000001111:
        _o_sv = 15'b111101010011000;
      13'b1101000010000:
        _o_sv = 15'b111101010011010;
      13'b1101000010001:
        _o_sv = 15'b111101010011011;
      13'b1101000010010:
        _o_sv = 15'b111101010011101;
      13'b1101000010011:
        _o_sv = 15'b111101010011111;
      13'b1101000010100:
        _o_sv = 15'b111101010100001;
      13'b1101000010101:
        _o_sv = 15'b111101010100011;
      13'b1101000010110:
        _o_sv = 15'b111101010100100;
      13'b1101000010111:
        _o_sv = 15'b111101010100110;
      13'b1101000011000:
        _o_sv = 15'b111101010101000;
      13'b1101000011001:
        _o_sv = 15'b111101010101010;
      13'b1101000011010:
        _o_sv = 15'b111101010101100;
      13'b1101000011011:
        _o_sv = 15'b111101010101101;
      13'b1101000011100:
        _o_sv = 15'b111101010101111;
      13'b1101000011101:
        _o_sv = 15'b111101010110001;
      13'b1101000011110:
        _o_sv = 15'b111101010110011;
      13'b1101000011111:
        _o_sv = 15'b111101010110101;
      13'b1101000100000:
        _o_sv = 15'b111101010110110;
      13'b1101000100001:
        _o_sv = 15'b111101010111000;
      13'b1101000100010:
        _o_sv = 15'b111101010111010;
      13'b1101000100011:
        _o_sv = 15'b111101010111100;
      13'b1101000100100:
        _o_sv = 15'b111101010111101;
      13'b1101000100101:
        _o_sv = 15'b111101010111111;
      13'b1101000100110:
        _o_sv = 15'b111101011000001;
      13'b1101000100111:
        _o_sv = 15'b111101011000011;
      13'b1101000101000:
        _o_sv = 15'b111101011000101;
      13'b1101000101001:
        _o_sv = 15'b111101011000110;
      13'b1101000101010:
        _o_sv = 15'b111101011001000;
      13'b1101000101011:
        _o_sv = 15'b111101011001010;
      13'b1101000101100:
        _o_sv = 15'b111101011001100;
      13'b1101000101101:
        _o_sv = 15'b111101011001101;
      13'b1101000101110:
        _o_sv = 15'b111101011001111;
      13'b1101000101111:
        _o_sv = 15'b111101011010001;
      13'b1101000110000:
        _o_sv = 15'b111101011010011;
      13'b1101000110001:
        _o_sv = 15'b111101011010101;
      13'b1101000110010:
        _o_sv = 15'b111101011010110;
      13'b1101000110011:
        _o_sv = 15'b111101011011000;
      13'b1101000110100:
        _o_sv = 15'b111101011011010;
      13'b1101000110101:
        _o_sv = 15'b111101011011100;
      13'b1101000110110:
        _o_sv = 15'b111101011011101;
      13'b1101000110111:
        _o_sv = 15'b111101011011111;
      13'b1101000111000:
        _o_sv = 15'b111101011100001;
      13'b1101000111001:
        _o_sv = 15'b111101011100011;
      13'b1101000111010:
        _o_sv = 15'b111101011100100;
      13'b1101000111011:
        _o_sv = 15'b111101011100110;
      13'b1101000111100:
        _o_sv = 15'b111101011101000;
      13'b1101000111101:
        _o_sv = 15'b111101011101010;
      13'b1101000111110:
        _o_sv = 15'b111101011101011;
      13'b1101000111111:
        _o_sv = 15'b111101011101101;
      13'b1101001000000:
        _o_sv = 15'b111101011101111;
      13'b1101001000001:
        _o_sv = 15'b111101011110001;
      13'b1101001000010:
        _o_sv = 15'b111101011110010;
      13'b1101001000011:
        _o_sv = 15'b111101011110100;
      13'b1101001000100:
        _o_sv = 15'b111101011110110;
      13'b1101001000101:
        _o_sv = 15'b111101011111000;
      13'b1101001000110:
        _o_sv = 15'b111101011111001;
      13'b1101001000111:
        _o_sv = 15'b111101011111011;
      13'b1101001001000:
        _o_sv = 15'b111101011111101;
      13'b1101001001001:
        _o_sv = 15'b111101011111111;
      13'b1101001001010:
        _o_sv = 15'b111101100000000;
      13'b1101001001011:
        _o_sv = 15'b111101100000010;
      13'b1101001001100:
        _o_sv = 15'b111101100000100;
      13'b1101001001101:
        _o_sv = 15'b111101100000110;
      13'b1101001001110:
        _o_sv = 15'b111101100000111;
      13'b1101001001111:
        _o_sv = 15'b111101100001001;
      13'b1101001010000:
        _o_sv = 15'b111101100001011;
      13'b1101001010001:
        _o_sv = 15'b111101100001100;
      13'b1101001010010:
        _o_sv = 15'b111101100001110;
      13'b1101001010011:
        _o_sv = 15'b111101100010000;
      13'b1101001010100:
        _o_sv = 15'b111101100010010;
      13'b1101001010101:
        _o_sv = 15'b111101100010011;
      13'b1101001010110:
        _o_sv = 15'b111101100010101;
      13'b1101001010111:
        _o_sv = 15'b111101100010111;
      13'b1101001011000:
        _o_sv = 15'b111101100011001;
      13'b1101001011001:
        _o_sv = 15'b111101100011010;
      13'b1101001011010:
        _o_sv = 15'b111101100011100;
      13'b1101001011011:
        _o_sv = 15'b111101100011110;
      13'b1101001011100:
        _o_sv = 15'b111101100011111;
      13'b1101001011101:
        _o_sv = 15'b111101100100001;
      13'b1101001011110:
        _o_sv = 15'b111101100100011;
      13'b1101001011111:
        _o_sv = 15'b111101100100101;
      13'b1101001100000:
        _o_sv = 15'b111101100100110;
      13'b1101001100001:
        _o_sv = 15'b111101100101000;
      13'b1101001100010:
        _o_sv = 15'b111101100101010;
      13'b1101001100011:
        _o_sv = 15'b111101100101011;
      13'b1101001100100:
        _o_sv = 15'b111101100101101;
      13'b1101001100101:
        _o_sv = 15'b111101100101111;
      13'b1101001100110:
        _o_sv = 15'b111101100110001;
      13'b1101001100111:
        _o_sv = 15'b111101100110010;
      13'b1101001101000:
        _o_sv = 15'b111101100110100;
      13'b1101001101001:
        _o_sv = 15'b111101100110110;
      13'b1101001101010:
        _o_sv = 15'b111101100110111;
      13'b1101001101011:
        _o_sv = 15'b111101100111001;
      13'b1101001101100:
        _o_sv = 15'b111101100111011;
      13'b1101001101101:
        _o_sv = 15'b111101100111100;
      13'b1101001101110:
        _o_sv = 15'b111101100111110;
      13'b1101001101111:
        _o_sv = 15'b111101101000000;
      13'b1101001110000:
        _o_sv = 15'b111101101000010;
      13'b1101001110001:
        _o_sv = 15'b111101101000011;
      13'b1101001110010:
        _o_sv = 15'b111101101000101;
      13'b1101001110011:
        _o_sv = 15'b111101101000111;
      13'b1101001110100:
        _o_sv = 15'b111101101001000;
      13'b1101001110101:
        _o_sv = 15'b111101101001010;
      13'b1101001110110:
        _o_sv = 15'b111101101001100;
      13'b1101001110111:
        _o_sv = 15'b111101101001101;
      13'b1101001111000:
        _o_sv = 15'b111101101001111;
      13'b1101001111001:
        _o_sv = 15'b111101101010001;
      13'b1101001111010:
        _o_sv = 15'b111101101010010;
      13'b1101001111011:
        _o_sv = 15'b111101101010100;
      13'b1101001111100:
        _o_sv = 15'b111101101010110;
      13'b1101001111101:
        _o_sv = 15'b111101101010111;
      13'b1101001111110:
        _o_sv = 15'b111101101011001;
      13'b1101001111111:
        _o_sv = 15'b111101101011011;
      13'b1101010000000:
        _o_sv = 15'b111101101011101;
      13'b1101010000001:
        _o_sv = 15'b111101101011110;
      13'b1101010000010:
        _o_sv = 15'b111101101100000;
      13'b1101010000011:
        _o_sv = 15'b111101101100010;
      13'b1101010000100:
        _o_sv = 15'b111101101100011;
      13'b1101010000101:
        _o_sv = 15'b111101101100101;
      13'b1101010000110:
        _o_sv = 15'b111101101100111;
      13'b1101010000111:
        _o_sv = 15'b111101101101000;
      13'b1101010001000:
        _o_sv = 15'b111101101101010;
      13'b1101010001001:
        _o_sv = 15'b111101101101100;
      13'b1101010001010:
        _o_sv = 15'b111101101101101;
      13'b1101010001011:
        _o_sv = 15'b111101101101111;
      13'b1101010001100:
        _o_sv = 15'b111101101110001;
      13'b1101010001101:
        _o_sv = 15'b111101101110010;
      13'b1101010001110:
        _o_sv = 15'b111101101110100;
      13'b1101010001111:
        _o_sv = 15'b111101101110110;
      13'b1101010010000:
        _o_sv = 15'b111101101110111;
      13'b1101010010001:
        _o_sv = 15'b111101101111001;
      13'b1101010010010:
        _o_sv = 15'b111101101111010;
      13'b1101010010011:
        _o_sv = 15'b111101101111100;
      13'b1101010010100:
        _o_sv = 15'b111101101111110;
      13'b1101010010101:
        _o_sv = 15'b111101101111111;
      13'b1101010010110:
        _o_sv = 15'b111101110000001;
      13'b1101010010111:
        _o_sv = 15'b111101110000011;
      13'b1101010011000:
        _o_sv = 15'b111101110000100;
      13'b1101010011001:
        _o_sv = 15'b111101110000110;
      13'b1101010011010:
        _o_sv = 15'b111101110001000;
      13'b1101010011011:
        _o_sv = 15'b111101110001001;
      13'b1101010011100:
        _o_sv = 15'b111101110001011;
      13'b1101010011101:
        _o_sv = 15'b111101110001101;
      13'b1101010011110:
        _o_sv = 15'b111101110001110;
      13'b1101010011111:
        _o_sv = 15'b111101110010000;
      13'b1101010100000:
        _o_sv = 15'b111101110010010;
      13'b1101010100001:
        _o_sv = 15'b111101110010011;
      13'b1101010100010:
        _o_sv = 15'b111101110010101;
      13'b1101010100011:
        _o_sv = 15'b111101110010110;
      13'b1101010100100:
        _o_sv = 15'b111101110011000;
      13'b1101010100101:
        _o_sv = 15'b111101110011010;
      13'b1101010100110:
        _o_sv = 15'b111101110011011;
      13'b1101010100111:
        _o_sv = 15'b111101110011101;
      13'b1101010101000:
        _o_sv = 15'b111101110011111;
      13'b1101010101001:
        _o_sv = 15'b111101110100000;
      13'b1101010101010:
        _o_sv = 15'b111101110100010;
      13'b1101010101011:
        _o_sv = 15'b111101110100011;
      13'b1101010101100:
        _o_sv = 15'b111101110100101;
      13'b1101010101101:
        _o_sv = 15'b111101110100111;
      13'b1101010101110:
        _o_sv = 15'b111101110101000;
      13'b1101010101111:
        _o_sv = 15'b111101110101010;
      13'b1101010110000:
        _o_sv = 15'b111101110101100;
      13'b1101010110001:
        _o_sv = 15'b111101110101101;
      13'b1101010110010:
        _o_sv = 15'b111101110101111;
      13'b1101010110011:
        _o_sv = 15'b111101110110000;
      13'b1101010110100:
        _o_sv = 15'b111101110110010;
      13'b1101010110101:
        _o_sv = 15'b111101110110100;
      13'b1101010110110:
        _o_sv = 15'b111101110110101;
      13'b1101010110111:
        _o_sv = 15'b111101110110111;
      13'b1101010111000:
        _o_sv = 15'b111101110111001;
      13'b1101010111001:
        _o_sv = 15'b111101110111010;
      13'b1101010111010:
        _o_sv = 15'b111101110111100;
      13'b1101010111011:
        _o_sv = 15'b111101110111101;
      13'b1101010111100:
        _o_sv = 15'b111101110111111;
      13'b1101010111101:
        _o_sv = 15'b111101111000001;
      13'b1101010111110:
        _o_sv = 15'b111101111000010;
      13'b1101010111111:
        _o_sv = 15'b111101111000100;
      13'b1101011000000:
        _o_sv = 15'b111101111000101;
      13'b1101011000001:
        _o_sv = 15'b111101111000111;
      13'b1101011000010:
        _o_sv = 15'b111101111001001;
      13'b1101011000011:
        _o_sv = 15'b111101111001010;
      13'b1101011000100:
        _o_sv = 15'b111101111001100;
      13'b1101011000101:
        _o_sv = 15'b111101111001101;
      13'b1101011000110:
        _o_sv = 15'b111101111001111;
      13'b1101011000111:
        _o_sv = 15'b111101111010001;
      13'b1101011001000:
        _o_sv = 15'b111101111010010;
      13'b1101011001001:
        _o_sv = 15'b111101111010100;
      13'b1101011001010:
        _o_sv = 15'b111101111010101;
      13'b1101011001011:
        _o_sv = 15'b111101111010111;
      13'b1101011001100:
        _o_sv = 15'b111101111011001;
      13'b1101011001101:
        _o_sv = 15'b111101111011010;
      13'b1101011001110:
        _o_sv = 15'b111101111011100;
      13'b1101011001111:
        _o_sv = 15'b111101111011101;
      13'b1101011010000:
        _o_sv = 15'b111101111011111;
      13'b1101011010001:
        _o_sv = 15'b111101111100000;
      13'b1101011010010:
        _o_sv = 15'b111101111100010;
      13'b1101011010011:
        _o_sv = 15'b111101111100100;
      13'b1101011010100:
        _o_sv = 15'b111101111100101;
      13'b1101011010101:
        _o_sv = 15'b111101111100111;
      13'b1101011010110:
        _o_sv = 15'b111101111101000;
      13'b1101011010111:
        _o_sv = 15'b111101111101010;
      13'b1101011011000:
        _o_sv = 15'b111101111101011;
      13'b1101011011001:
        _o_sv = 15'b111101111101101;
      13'b1101011011010:
        _o_sv = 15'b111101111101111;
      13'b1101011011011:
        _o_sv = 15'b111101111110000;
      13'b1101011011100:
        _o_sv = 15'b111101111110010;
      13'b1101011011101:
        _o_sv = 15'b111101111110011;
      13'b1101011011110:
        _o_sv = 15'b111101111110101;
      13'b1101011011111:
        _o_sv = 15'b111101111110110;
      13'b1101011100000:
        _o_sv = 15'b111101111111000;
      13'b1101011100001:
        _o_sv = 15'b111101111111010;
      13'b1101011100010:
        _o_sv = 15'b111101111111011;
      13'b1101011100011:
        _o_sv = 15'b111101111111101;
      13'b1101011100100:
        _o_sv = 15'b111101111111110;
      13'b1101011100101:
        _o_sv = 15'b111110000000000;
      13'b1101011100110:
        _o_sv = 15'b111110000000001;
      13'b1101011100111:
        _o_sv = 15'b111110000000011;
      13'b1101011101000:
        _o_sv = 15'b111110000000101;
      13'b1101011101001:
        _o_sv = 15'b111110000000110;
      13'b1101011101010:
        _o_sv = 15'b111110000001000;
      13'b1101011101011:
        _o_sv = 15'b111110000001001;
      13'b1101011101100:
        _o_sv = 15'b111110000001011;
      13'b1101011101101:
        _o_sv = 15'b111110000001100;
      13'b1101011101110:
        _o_sv = 15'b111110000001110;
      13'b1101011101111:
        _o_sv = 15'b111110000001111;
      13'b1101011110000:
        _o_sv = 15'b111110000010001;
      13'b1101011110001:
        _o_sv = 15'b111110000010010;
      13'b1101011110010:
        _o_sv = 15'b111110000010100;
      13'b1101011110011:
        _o_sv = 15'b111110000010110;
      13'b1101011110100:
        _o_sv = 15'b111110000010111;
      13'b1101011110101:
        _o_sv = 15'b111110000011001;
      13'b1101011110110:
        _o_sv = 15'b111110000011010;
      13'b1101011110111:
        _o_sv = 15'b111110000011100;
      13'b1101011111000:
        _o_sv = 15'b111110000011101;
      13'b1101011111001:
        _o_sv = 15'b111110000011111;
      13'b1101011111010:
        _o_sv = 15'b111110000100000;
      13'b1101011111011:
        _o_sv = 15'b111110000100010;
      13'b1101011111100:
        _o_sv = 15'b111110000100011;
      13'b1101011111101:
        _o_sv = 15'b111110000100101;
      13'b1101011111110:
        _o_sv = 15'b111110000100110;
      13'b1101011111111:
        _o_sv = 15'b111110000101000;
      13'b1101100000000:
        _o_sv = 15'b111110000101001;
      13'b1101100000001:
        _o_sv = 15'b111110000101011;
      13'b1101100000010:
        _o_sv = 15'b111110000101101;
      13'b1101100000011:
        _o_sv = 15'b111110000101110;
      13'b1101100000100:
        _o_sv = 15'b111110000110000;
      13'b1101100000101:
        _o_sv = 15'b111110000110001;
      13'b1101100000110:
        _o_sv = 15'b111110000110011;
      13'b1101100000111:
        _o_sv = 15'b111110000110100;
      13'b1101100001000:
        _o_sv = 15'b111110000110110;
      13'b1101100001001:
        _o_sv = 15'b111110000110111;
      13'b1101100001010:
        _o_sv = 15'b111110000111001;
      13'b1101100001011:
        _o_sv = 15'b111110000111010;
      13'b1101100001100:
        _o_sv = 15'b111110000111100;
      13'b1101100001101:
        _o_sv = 15'b111110000111101;
      13'b1101100001110:
        _o_sv = 15'b111110000111111;
      13'b1101100001111:
        _o_sv = 15'b111110001000000;
      13'b1101100010000:
        _o_sv = 15'b111110001000010;
      13'b1101100010001:
        _o_sv = 15'b111110001000011;
      13'b1101100010010:
        _o_sv = 15'b111110001000101;
      13'b1101100010011:
        _o_sv = 15'b111110001000110;
      13'b1101100010100:
        _o_sv = 15'b111110001001000;
      13'b1101100010101:
        _o_sv = 15'b111110001001001;
      13'b1101100010110:
        _o_sv = 15'b111110001001011;
      13'b1101100010111:
        _o_sv = 15'b111110001001100;
      13'b1101100011000:
        _o_sv = 15'b111110001001110;
      13'b1101100011001:
        _o_sv = 15'b111110001001111;
      13'b1101100011010:
        _o_sv = 15'b111110001010001;
      13'b1101100011011:
        _o_sv = 15'b111110001010010;
      13'b1101100011100:
        _o_sv = 15'b111110001010100;
      13'b1101100011101:
        _o_sv = 15'b111110001010101;
      13'b1101100011110:
        _o_sv = 15'b111110001010111;
      13'b1101100011111:
        _o_sv = 15'b111110001011000;
      13'b1101100100000:
        _o_sv = 15'b111110001011010;
      13'b1101100100001:
        _o_sv = 15'b111110001011011;
      13'b1101100100010:
        _o_sv = 15'b111110001011101;
      13'b1101100100011:
        _o_sv = 15'b111110001011110;
      13'b1101100100100:
        _o_sv = 15'b111110001100000;
      13'b1101100100101:
        _o_sv = 15'b111110001100001;
      13'b1101100100110:
        _o_sv = 15'b111110001100011;
      13'b1101100100111:
        _o_sv = 15'b111110001100100;
      13'b1101100101000:
        _o_sv = 15'b111110001100110;
      13'b1101100101001:
        _o_sv = 15'b111110001100111;
      13'b1101100101010:
        _o_sv = 15'b111110001101001;
      13'b1101100101011:
        _o_sv = 15'b111110001101010;
      13'b1101100101100:
        _o_sv = 15'b111110001101100;
      13'b1101100101101:
        _o_sv = 15'b111110001101101;
      13'b1101100101110:
        _o_sv = 15'b111110001101110;
      13'b1101100101111:
        _o_sv = 15'b111110001110000;
      13'b1101100110000:
        _o_sv = 15'b111110001110001;
      13'b1101100110001:
        _o_sv = 15'b111110001110011;
      13'b1101100110010:
        _o_sv = 15'b111110001110100;
      13'b1101100110011:
        _o_sv = 15'b111110001110110;
      13'b1101100110100:
        _o_sv = 15'b111110001110111;
      13'b1101100110101:
        _o_sv = 15'b111110001111001;
      13'b1101100110110:
        _o_sv = 15'b111110001111010;
      13'b1101100110111:
        _o_sv = 15'b111110001111100;
      13'b1101100111000:
        _o_sv = 15'b111110001111101;
      13'b1101100111001:
        _o_sv = 15'b111110001111111;
      13'b1101100111010:
        _o_sv = 15'b111110010000000;
      13'b1101100111011:
        _o_sv = 15'b111110010000010;
      13'b1101100111100:
        _o_sv = 15'b111110010000011;
      13'b1101100111101:
        _o_sv = 15'b111110010000100;
      13'b1101100111110:
        _o_sv = 15'b111110010000110;
      13'b1101100111111:
        _o_sv = 15'b111110010000111;
      13'b1101101000000:
        _o_sv = 15'b111110010001001;
      13'b1101101000001:
        _o_sv = 15'b111110010001010;
      13'b1101101000010:
        _o_sv = 15'b111110010001100;
      13'b1101101000011:
        _o_sv = 15'b111110010001101;
      13'b1101101000100:
        _o_sv = 15'b111110010001111;
      13'b1101101000101:
        _o_sv = 15'b111110010010000;
      13'b1101101000110:
        _o_sv = 15'b111110010010001;
      13'b1101101000111:
        _o_sv = 15'b111110010010011;
      13'b1101101001000:
        _o_sv = 15'b111110010010100;
      13'b1101101001001:
        _o_sv = 15'b111110010010110;
      13'b1101101001010:
        _o_sv = 15'b111110010010111;
      13'b1101101001011:
        _o_sv = 15'b111110010011001;
      13'b1101101001100:
        _o_sv = 15'b111110010011010;
      13'b1101101001101:
        _o_sv = 15'b111110010011100;
      13'b1101101001110:
        _o_sv = 15'b111110010011101;
      13'b1101101001111:
        _o_sv = 15'b111110010011110;
      13'b1101101010000:
        _o_sv = 15'b111110010100000;
      13'b1101101010001:
        _o_sv = 15'b111110010100001;
      13'b1101101010010:
        _o_sv = 15'b111110010100011;
      13'b1101101010011:
        _o_sv = 15'b111110010100100;
      13'b1101101010100:
        _o_sv = 15'b111110010100110;
      13'b1101101010101:
        _o_sv = 15'b111110010100111;
      13'b1101101010110:
        _o_sv = 15'b111110010101000;
      13'b1101101010111:
        _o_sv = 15'b111110010101010;
      13'b1101101011000:
        _o_sv = 15'b111110010101011;
      13'b1101101011001:
        _o_sv = 15'b111110010101101;
      13'b1101101011010:
        _o_sv = 15'b111110010101110;
      13'b1101101011011:
        _o_sv = 15'b111110010110000;
      13'b1101101011100:
        _o_sv = 15'b111110010110001;
      13'b1101101011101:
        _o_sv = 15'b111110010110010;
      13'b1101101011110:
        _o_sv = 15'b111110010110100;
      13'b1101101011111:
        _o_sv = 15'b111110010110101;
      13'b1101101100000:
        _o_sv = 15'b111110010110111;
      13'b1101101100001:
        _o_sv = 15'b111110010111000;
      13'b1101101100010:
        _o_sv = 15'b111110010111001;
      13'b1101101100011:
        _o_sv = 15'b111110010111011;
      13'b1101101100100:
        _o_sv = 15'b111110010111100;
      13'b1101101100101:
        _o_sv = 15'b111110010111110;
      13'b1101101100110:
        _o_sv = 15'b111110010111111;
      13'b1101101100111:
        _o_sv = 15'b111110011000001;
      13'b1101101101000:
        _o_sv = 15'b111110011000010;
      13'b1101101101001:
        _o_sv = 15'b111110011000011;
      13'b1101101101010:
        _o_sv = 15'b111110011000101;
      13'b1101101101011:
        _o_sv = 15'b111110011000110;
      13'b1101101101100:
        _o_sv = 15'b111110011001000;
      13'b1101101101101:
        _o_sv = 15'b111110011001001;
      13'b1101101101110:
        _o_sv = 15'b111110011001010;
      13'b1101101101111:
        _o_sv = 15'b111110011001100;
      13'b1101101110000:
        _o_sv = 15'b111110011001101;
      13'b1101101110001:
        _o_sv = 15'b111110011001111;
      13'b1101101110010:
        _o_sv = 15'b111110011010000;
      13'b1101101110011:
        _o_sv = 15'b111110011010001;
      13'b1101101110100:
        _o_sv = 15'b111110011010011;
      13'b1101101110101:
        _o_sv = 15'b111110011010100;
      13'b1101101110110:
        _o_sv = 15'b111110011010101;
      13'b1101101110111:
        _o_sv = 15'b111110011010111;
      13'b1101101111000:
        _o_sv = 15'b111110011011000;
      13'b1101101111001:
        _o_sv = 15'b111110011011010;
      13'b1101101111010:
        _o_sv = 15'b111110011011011;
      13'b1101101111011:
        _o_sv = 15'b111110011011100;
      13'b1101101111100:
        _o_sv = 15'b111110011011110;
      13'b1101101111101:
        _o_sv = 15'b111110011011111;
      13'b1101101111110:
        _o_sv = 15'b111110011100001;
      13'b1101101111111:
        _o_sv = 15'b111110011100010;
      13'b1101110000000:
        _o_sv = 15'b111110011100011;
      13'b1101110000001:
        _o_sv = 15'b111110011100101;
      13'b1101110000010:
        _o_sv = 15'b111110011100110;
      13'b1101110000011:
        _o_sv = 15'b111110011100111;
      13'b1101110000100:
        _o_sv = 15'b111110011101001;
      13'b1101110000101:
        _o_sv = 15'b111110011101010;
      13'b1101110000110:
        _o_sv = 15'b111110011101100;
      13'b1101110000111:
        _o_sv = 15'b111110011101101;
      13'b1101110001000:
        _o_sv = 15'b111110011101110;
      13'b1101110001001:
        _o_sv = 15'b111110011110000;
      13'b1101110001010:
        _o_sv = 15'b111110011110001;
      13'b1101110001011:
        _o_sv = 15'b111110011110010;
      13'b1101110001100:
        _o_sv = 15'b111110011110100;
      13'b1101110001101:
        _o_sv = 15'b111110011110101;
      13'b1101110001110:
        _o_sv = 15'b111110011110110;
      13'b1101110001111:
        _o_sv = 15'b111110011111000;
      13'b1101110010000:
        _o_sv = 15'b111110011111001;
      13'b1101110010001:
        _o_sv = 15'b111110011111011;
      13'b1101110010010:
        _o_sv = 15'b111110011111100;
      13'b1101110010011:
        _o_sv = 15'b111110011111101;
      13'b1101110010100:
        _o_sv = 15'b111110011111111;
      13'b1101110010101:
        _o_sv = 15'b111110100000000;
      13'b1101110010110:
        _o_sv = 15'b111110100000001;
      13'b1101110010111:
        _o_sv = 15'b111110100000011;
      13'b1101110011000:
        _o_sv = 15'b111110100000100;
      13'b1101110011001:
        _o_sv = 15'b111110100000101;
      13'b1101110011010:
        _o_sv = 15'b111110100000111;
      13'b1101110011011:
        _o_sv = 15'b111110100001000;
      13'b1101110011100:
        _o_sv = 15'b111110100001001;
      13'b1101110011101:
        _o_sv = 15'b111110100001011;
      13'b1101110011110:
        _o_sv = 15'b111110100001100;
      13'b1101110011111:
        _o_sv = 15'b111110100001101;
      13'b1101110100000:
        _o_sv = 15'b111110100001111;
      13'b1101110100001:
        _o_sv = 15'b111110100010000;
      13'b1101110100010:
        _o_sv = 15'b111110100010001;
      13'b1101110100011:
        _o_sv = 15'b111110100010011;
      13'b1101110100100:
        _o_sv = 15'b111110100010100;
      13'b1101110100101:
        _o_sv = 15'b111110100010101;
      13'b1101110100110:
        _o_sv = 15'b111110100010111;
      13'b1101110100111:
        _o_sv = 15'b111110100011000;
      13'b1101110101000:
        _o_sv = 15'b111110100011001;
      13'b1101110101001:
        _o_sv = 15'b111110100011011;
      13'b1101110101010:
        _o_sv = 15'b111110100011100;
      13'b1101110101011:
        _o_sv = 15'b111110100011101;
      13'b1101110101100:
        _o_sv = 15'b111110100011111;
      13'b1101110101101:
        _o_sv = 15'b111110100100000;
      13'b1101110101110:
        _o_sv = 15'b111110100100001;
      13'b1101110101111:
        _o_sv = 15'b111110100100011;
      13'b1101110110000:
        _o_sv = 15'b111110100100100;
      13'b1101110110001:
        _o_sv = 15'b111110100100101;
      13'b1101110110010:
        _o_sv = 15'b111110100100111;
      13'b1101110110011:
        _o_sv = 15'b111110100101000;
      13'b1101110110100:
        _o_sv = 15'b111110100101001;
      13'b1101110110101:
        _o_sv = 15'b111110100101011;
      13'b1101110110110:
        _o_sv = 15'b111110100101100;
      13'b1101110110111:
        _o_sv = 15'b111110100101101;
      13'b1101110111000:
        _o_sv = 15'b111110100101111;
      13'b1101110111001:
        _o_sv = 15'b111110100110000;
      13'b1101110111010:
        _o_sv = 15'b111110100110001;
      13'b1101110111011:
        _o_sv = 15'b111110100110010;
      13'b1101110111100:
        _o_sv = 15'b111110100110100;
      13'b1101110111101:
        _o_sv = 15'b111110100110101;
      13'b1101110111110:
        _o_sv = 15'b111110100110110;
      13'b1101110111111:
        _o_sv = 15'b111110100111000;
      13'b1101111000000:
        _o_sv = 15'b111110100111001;
      13'b1101111000001:
        _o_sv = 15'b111110100111010;
      13'b1101111000010:
        _o_sv = 15'b111110100111100;
      13'b1101111000011:
        _o_sv = 15'b111110100111101;
      13'b1101111000100:
        _o_sv = 15'b111110100111110;
      13'b1101111000101:
        _o_sv = 15'b111110100111111;
      13'b1101111000110:
        _o_sv = 15'b111110101000001;
      13'b1101111000111:
        _o_sv = 15'b111110101000010;
      13'b1101111001000:
        _o_sv = 15'b111110101000011;
      13'b1101111001001:
        _o_sv = 15'b111110101000101;
      13'b1101111001010:
        _o_sv = 15'b111110101000110;
      13'b1101111001011:
        _o_sv = 15'b111110101000111;
      13'b1101111001100:
        _o_sv = 15'b111110101001001;
      13'b1101111001101:
        _o_sv = 15'b111110101001010;
      13'b1101111001110:
        _o_sv = 15'b111110101001011;
      13'b1101111001111:
        _o_sv = 15'b111110101001100;
      13'b1101111010000:
        _o_sv = 15'b111110101001110;
      13'b1101111010001:
        _o_sv = 15'b111110101001111;
      13'b1101111010010:
        _o_sv = 15'b111110101010000;
      13'b1101111010011:
        _o_sv = 15'b111110101010010;
      13'b1101111010100:
        _o_sv = 15'b111110101010011;
      13'b1101111010101:
        _o_sv = 15'b111110101010100;
      13'b1101111010110:
        _o_sv = 15'b111110101010101;
      13'b1101111010111:
        _o_sv = 15'b111110101010111;
      13'b1101111011000:
        _o_sv = 15'b111110101011000;
      13'b1101111011001:
        _o_sv = 15'b111110101011001;
      13'b1101111011010:
        _o_sv = 15'b111110101011010;
      13'b1101111011011:
        _o_sv = 15'b111110101011100;
      13'b1101111011100:
        _o_sv = 15'b111110101011101;
      13'b1101111011101:
        _o_sv = 15'b111110101011110;
      13'b1101111011110:
        _o_sv = 15'b111110101100000;
      13'b1101111011111:
        _o_sv = 15'b111110101100001;
      13'b1101111100000:
        _o_sv = 15'b111110101100010;
      13'b1101111100001:
        _o_sv = 15'b111110101100011;
      13'b1101111100010:
        _o_sv = 15'b111110101100101;
      13'b1101111100011:
        _o_sv = 15'b111110101100110;
      13'b1101111100100:
        _o_sv = 15'b111110101100111;
      13'b1101111100101:
        _o_sv = 15'b111110101101000;
      13'b1101111100110:
        _o_sv = 15'b111110101101010;
      13'b1101111100111:
        _o_sv = 15'b111110101101011;
      13'b1101111101000:
        _o_sv = 15'b111110101101100;
      13'b1101111101001:
        _o_sv = 15'b111110101101101;
      13'b1101111101010:
        _o_sv = 15'b111110101101111;
      13'b1101111101011:
        _o_sv = 15'b111110101110000;
      13'b1101111101100:
        _o_sv = 15'b111110101110001;
      13'b1101111101101:
        _o_sv = 15'b111110101110010;
      13'b1101111101110:
        _o_sv = 15'b111110101110100;
      13'b1101111101111:
        _o_sv = 15'b111110101110101;
      13'b1101111110000:
        _o_sv = 15'b111110101110110;
      13'b1101111110001:
        _o_sv = 15'b111110101110111;
      13'b1101111110010:
        _o_sv = 15'b111110101111001;
      13'b1101111110011:
        _o_sv = 15'b111110101111010;
      13'b1101111110100:
        _o_sv = 15'b111110101111011;
      13'b1101111110101:
        _o_sv = 15'b111110101111100;
      13'b1101111110110:
        _o_sv = 15'b111110101111110;
      13'b1101111110111:
        _o_sv = 15'b111110101111111;
      13'b1101111111000:
        _o_sv = 15'b111110110000000;
      13'b1101111111001:
        _o_sv = 15'b111110110000001;
      13'b1101111111010:
        _o_sv = 15'b111110110000010;
      13'b1101111111011:
        _o_sv = 15'b111110110000100;
      13'b1101111111100:
        _o_sv = 15'b111110110000101;
      13'b1101111111101:
        _o_sv = 15'b111110110000110;
      13'b1101111111110:
        _o_sv = 15'b111110110000111;
      13'b1101111111111:
        _o_sv = 15'b111110110001001;
      13'b1110000000000:
        _o_sv = 15'b111110110001010;
      13'b1110000000001:
        _o_sv = 15'b111110110001011;
      13'b1110000000010:
        _o_sv = 15'b111110110001100;
      13'b1110000000011:
        _o_sv = 15'b111110110001110;
      13'b1110000000100:
        _o_sv = 15'b111110110001111;
      13'b1110000000101:
        _o_sv = 15'b111110110010000;
      13'b1110000000110:
        _o_sv = 15'b111110110010001;
      13'b1110000000111:
        _o_sv = 15'b111110110010010;
      13'b1110000001000:
        _o_sv = 15'b111110110010100;
      13'b1110000001001:
        _o_sv = 15'b111110110010101;
      13'b1110000001010:
        _o_sv = 15'b111110110010110;
      13'b1110000001011:
        _o_sv = 15'b111110110010111;
      13'b1110000001100:
        _o_sv = 15'b111110110011000;
      13'b1110000001101:
        _o_sv = 15'b111110110011010;
      13'b1110000001110:
        _o_sv = 15'b111110110011011;
      13'b1110000001111:
        _o_sv = 15'b111110110011100;
      13'b1110000010000:
        _o_sv = 15'b111110110011101;
      13'b1110000010001:
        _o_sv = 15'b111110110011111;
      13'b1110000010010:
        _o_sv = 15'b111110110100000;
      13'b1110000010011:
        _o_sv = 15'b111110110100001;
      13'b1110000010100:
        _o_sv = 15'b111110110100010;
      13'b1110000010101:
        _o_sv = 15'b111110110100011;
      13'b1110000010110:
        _o_sv = 15'b111110110100101;
      13'b1110000010111:
        _o_sv = 15'b111110110100110;
      13'b1110000011000:
        _o_sv = 15'b111110110100111;
      13'b1110000011001:
        _o_sv = 15'b111110110101000;
      13'b1110000011010:
        _o_sv = 15'b111110110101001;
      13'b1110000011011:
        _o_sv = 15'b111110110101011;
      13'b1110000011100:
        _o_sv = 15'b111110110101100;
      13'b1110000011101:
        _o_sv = 15'b111110110101101;
      13'b1110000011110:
        _o_sv = 15'b111110110101110;
      13'b1110000011111:
        _o_sv = 15'b111110110101111;
      13'b1110000100000:
        _o_sv = 15'b111110110110000;
      13'b1110000100001:
        _o_sv = 15'b111110110110010;
      13'b1110000100010:
        _o_sv = 15'b111110110110011;
      13'b1110000100011:
        _o_sv = 15'b111110110110100;
      13'b1110000100100:
        _o_sv = 15'b111110110110101;
      13'b1110000100101:
        _o_sv = 15'b111110110110110;
      13'b1110000100110:
        _o_sv = 15'b111110110111000;
      13'b1110000100111:
        _o_sv = 15'b111110110111001;
      13'b1110000101000:
        _o_sv = 15'b111110110111010;
      13'b1110000101001:
        _o_sv = 15'b111110110111011;
      13'b1110000101010:
        _o_sv = 15'b111110110111100;
      13'b1110000101011:
        _o_sv = 15'b111110110111101;
      13'b1110000101100:
        _o_sv = 15'b111110110111111;
      13'b1110000101101:
        _o_sv = 15'b111110111000000;
      13'b1110000101110:
        _o_sv = 15'b111110111000001;
      13'b1110000101111:
        _o_sv = 15'b111110111000010;
      13'b1110000110000:
        _o_sv = 15'b111110111000011;
      13'b1110000110001:
        _o_sv = 15'b111110111000101;
      13'b1110000110010:
        _o_sv = 15'b111110111000110;
      13'b1110000110011:
        _o_sv = 15'b111110111000111;
      13'b1110000110100:
        _o_sv = 15'b111110111001000;
      13'b1110000110101:
        _o_sv = 15'b111110111001001;
      13'b1110000110110:
        _o_sv = 15'b111110111001010;
      13'b1110000110111:
        _o_sv = 15'b111110111001100;
      13'b1110000111000:
        _o_sv = 15'b111110111001101;
      13'b1110000111001:
        _o_sv = 15'b111110111001110;
      13'b1110000111010:
        _o_sv = 15'b111110111001111;
      13'b1110000111011:
        _o_sv = 15'b111110111010000;
      13'b1110000111100:
        _o_sv = 15'b111110111010001;
      13'b1110000111101:
        _o_sv = 15'b111110111010010;
      13'b1110000111110:
        _o_sv = 15'b111110111010100;
      13'b1110000111111:
        _o_sv = 15'b111110111010101;
      13'b1110001000000:
        _o_sv = 15'b111110111010110;
      13'b1110001000001:
        _o_sv = 15'b111110111010111;
      13'b1110001000010:
        _o_sv = 15'b111110111011000;
      13'b1110001000011:
        _o_sv = 15'b111110111011001;
      13'b1110001000100:
        _o_sv = 15'b111110111011010;
      13'b1110001000101:
        _o_sv = 15'b111110111011100;
      13'b1110001000110:
        _o_sv = 15'b111110111011101;
      13'b1110001000111:
        _o_sv = 15'b111110111011110;
      13'b1110001001000:
        _o_sv = 15'b111110111011111;
      13'b1110001001001:
        _o_sv = 15'b111110111100000;
      13'b1110001001010:
        _o_sv = 15'b111110111100001;
      13'b1110001001011:
        _o_sv = 15'b111110111100010;
      13'b1110001001100:
        _o_sv = 15'b111110111100100;
      13'b1110001001101:
        _o_sv = 15'b111110111100101;
      13'b1110001001110:
        _o_sv = 15'b111110111100110;
      13'b1110001001111:
        _o_sv = 15'b111110111100111;
      13'b1110001010000:
        _o_sv = 15'b111110111101000;
      13'b1110001010001:
        _o_sv = 15'b111110111101001;
      13'b1110001010010:
        _o_sv = 15'b111110111101010;
      13'b1110001010011:
        _o_sv = 15'b111110111101100;
      13'b1110001010100:
        _o_sv = 15'b111110111101101;
      13'b1110001010101:
        _o_sv = 15'b111110111101110;
      13'b1110001010110:
        _o_sv = 15'b111110111101111;
      13'b1110001010111:
        _o_sv = 15'b111110111110000;
      13'b1110001011000:
        _o_sv = 15'b111110111110001;
      13'b1110001011001:
        _o_sv = 15'b111110111110010;
      13'b1110001011010:
        _o_sv = 15'b111110111110011;
      13'b1110001011011:
        _o_sv = 15'b111110111110101;
      13'b1110001011100:
        _o_sv = 15'b111110111110110;
      13'b1110001011101:
        _o_sv = 15'b111110111110111;
      13'b1110001011110:
        _o_sv = 15'b111110111111000;
      13'b1110001011111:
        _o_sv = 15'b111110111111001;
      13'b1110001100000:
        _o_sv = 15'b111110111111010;
      13'b1110001100001:
        _o_sv = 15'b111110111111011;
      13'b1110001100010:
        _o_sv = 15'b111110111111100;
      13'b1110001100011:
        _o_sv = 15'b111110111111101;
      13'b1110001100100:
        _o_sv = 15'b111110111111111;
      13'b1110001100101:
        _o_sv = 15'b111111000000000;
      13'b1110001100110:
        _o_sv = 15'b111111000000001;
      13'b1110001100111:
        _o_sv = 15'b111111000000010;
      13'b1110001101000:
        _o_sv = 15'b111111000000011;
      13'b1110001101001:
        _o_sv = 15'b111111000000100;
      13'b1110001101010:
        _o_sv = 15'b111111000000101;
      13'b1110001101011:
        _o_sv = 15'b111111000000110;
      13'b1110001101100:
        _o_sv = 15'b111111000000111;
      13'b1110001101101:
        _o_sv = 15'b111111000001000;
      13'b1110001101110:
        _o_sv = 15'b111111000001010;
      13'b1110001101111:
        _o_sv = 15'b111111000001011;
      13'b1110001110000:
        _o_sv = 15'b111111000001100;
      13'b1110001110001:
        _o_sv = 15'b111111000001101;
      13'b1110001110010:
        _o_sv = 15'b111111000001110;
      13'b1110001110011:
        _o_sv = 15'b111111000001111;
      13'b1110001110100:
        _o_sv = 15'b111111000010000;
      13'b1110001110101:
        _o_sv = 15'b111111000010001;
      13'b1110001110110:
        _o_sv = 15'b111111000010010;
      13'b1110001110111:
        _o_sv = 15'b111111000010011;
      13'b1110001111000:
        _o_sv = 15'b111111000010100;
      13'b1110001111001:
        _o_sv = 15'b111111000010110;
      13'b1110001111010:
        _o_sv = 15'b111111000010111;
      13'b1110001111011:
        _o_sv = 15'b111111000011000;
      13'b1110001111100:
        _o_sv = 15'b111111000011001;
      13'b1110001111101:
        _o_sv = 15'b111111000011010;
      13'b1110001111110:
        _o_sv = 15'b111111000011011;
      13'b1110001111111:
        _o_sv = 15'b111111000011100;
      13'b1110010000000:
        _o_sv = 15'b111111000011101;
      13'b1110010000001:
        _o_sv = 15'b111111000011110;
      13'b1110010000010:
        _o_sv = 15'b111111000011111;
      13'b1110010000011:
        _o_sv = 15'b111111000100000;
      13'b1110010000100:
        _o_sv = 15'b111111000100001;
      13'b1110010000101:
        _o_sv = 15'b111111000100010;
      13'b1110010000110:
        _o_sv = 15'b111111000100100;
      13'b1110010000111:
        _o_sv = 15'b111111000100101;
      13'b1110010001000:
        _o_sv = 15'b111111000100110;
      13'b1110010001001:
        _o_sv = 15'b111111000100111;
      13'b1110010001010:
        _o_sv = 15'b111111000101000;
      13'b1110010001011:
        _o_sv = 15'b111111000101001;
      13'b1110010001100:
        _o_sv = 15'b111111000101010;
      13'b1110010001101:
        _o_sv = 15'b111111000101011;
      13'b1110010001110:
        _o_sv = 15'b111111000101100;
      13'b1110010001111:
        _o_sv = 15'b111111000101101;
      13'b1110010010000:
        _o_sv = 15'b111111000101110;
      13'b1110010010001:
        _o_sv = 15'b111111000101111;
      13'b1110010010010:
        _o_sv = 15'b111111000110000;
      13'b1110010010011:
        _o_sv = 15'b111111000110001;
      13'b1110010010100:
        _o_sv = 15'b111111000110010;
      13'b1110010010101:
        _o_sv = 15'b111111000110011;
      13'b1110010010110:
        _o_sv = 15'b111111000110100;
      13'b1110010010111:
        _o_sv = 15'b111111000110101;
      13'b1110010011000:
        _o_sv = 15'b111111000110111;
      13'b1110010011001:
        _o_sv = 15'b111111000111000;
      13'b1110010011010:
        _o_sv = 15'b111111000111001;
      13'b1110010011011:
        _o_sv = 15'b111111000111010;
      13'b1110010011100:
        _o_sv = 15'b111111000111011;
      13'b1110010011101:
        _o_sv = 15'b111111000111100;
      13'b1110010011110:
        _o_sv = 15'b111111000111101;
      13'b1110010011111:
        _o_sv = 15'b111111000111110;
      13'b1110010100000:
        _o_sv = 15'b111111000111111;
      13'b1110010100001:
        _o_sv = 15'b111111001000000;
      13'b1110010100010:
        _o_sv = 15'b111111001000001;
      13'b1110010100011:
        _o_sv = 15'b111111001000010;
      13'b1110010100100:
        _o_sv = 15'b111111001000011;
      13'b1110010100101:
        _o_sv = 15'b111111001000100;
      13'b1110010100110:
        _o_sv = 15'b111111001000101;
      13'b1110010100111:
        _o_sv = 15'b111111001000110;
      13'b1110010101000:
        _o_sv = 15'b111111001000111;
      13'b1110010101001:
        _o_sv = 15'b111111001001000;
      13'b1110010101010:
        _o_sv = 15'b111111001001001;
      13'b1110010101011:
        _o_sv = 15'b111111001001010;
      13'b1110010101100:
        _o_sv = 15'b111111001001011;
      13'b1110010101101:
        _o_sv = 15'b111111001001100;
      13'b1110010101110:
        _o_sv = 15'b111111001001101;
      13'b1110010101111:
        _o_sv = 15'b111111001001110;
      13'b1110010110000:
        _o_sv = 15'b111111001001111;
      13'b1110010110001:
        _o_sv = 15'b111111001010000;
      13'b1110010110010:
        _o_sv = 15'b111111001010001;
      13'b1110010110011:
        _o_sv = 15'b111111001010010;
      13'b1110010110100:
        _o_sv = 15'b111111001010011;
      13'b1110010110101:
        _o_sv = 15'b111111001010100;
      13'b1110010110110:
        _o_sv = 15'b111111001010101;
      13'b1110010110111:
        _o_sv = 15'b111111001010110;
      13'b1110010111000:
        _o_sv = 15'b111111001010111;
      13'b1110010111001:
        _o_sv = 15'b111111001011000;
      13'b1110010111010:
        _o_sv = 15'b111111001011001;
      13'b1110010111011:
        _o_sv = 15'b111111001011010;
      13'b1110010111100:
        _o_sv = 15'b111111001011011;
      13'b1110010111101:
        _o_sv = 15'b111111001011100;
      13'b1110010111110:
        _o_sv = 15'b111111001011101;
      13'b1110010111111:
        _o_sv = 15'b111111001011110;
      13'b1110011000000:
        _o_sv = 15'b111111001011111;
      13'b1110011000001:
        _o_sv = 15'b111111001100000;
      13'b1110011000010:
        _o_sv = 15'b111111001100001;
      13'b1110011000011:
        _o_sv = 15'b111111001100010;
      13'b1110011000100:
        _o_sv = 15'b111111001100011;
      13'b1110011000101:
        _o_sv = 15'b111111001100100;
      13'b1110011000110:
        _o_sv = 15'b111111001100101;
      13'b1110011000111:
        _o_sv = 15'b111111001100110;
      13'b1110011001000:
        _o_sv = 15'b111111001100111;
      13'b1110011001001:
        _o_sv = 15'b111111001101000;
      13'b1110011001010:
        _o_sv = 15'b111111001101001;
      13'b1110011001011:
        _o_sv = 15'b111111001101010;
      13'b1110011001100:
        _o_sv = 15'b111111001101011;
      13'b1110011001101:
        _o_sv = 15'b111111001101100;
      13'b1110011001110:
        _o_sv = 15'b111111001101101;
      13'b1110011001111:
        _o_sv = 15'b111111001101110;
      13'b1110011010000:
        _o_sv = 15'b111111001101111;
      13'b1110011010001:
        _o_sv = 15'b111111001110000;
      13'b1110011010010:
        _o_sv = 15'b111111001110001;
      13'b1110011010011:
        _o_sv = 15'b111111001110010;
      13'b1110011010100:
        _o_sv = 15'b111111001110011;
      13'b1110011010101:
        _o_sv = 15'b111111001110100;
      13'b1110011010110:
        _o_sv = 15'b111111001110101;
      13'b1110011010111:
        _o_sv = 15'b111111001110110;
      13'b1110011011000:
        _o_sv = 15'b111111001110111;
      13'b1110011011001:
        _o_sv = 15'b111111001111000;
      13'b1110011011010:
        _o_sv = 15'b111111001111001;
      13'b1110011011011:
        _o_sv = 15'b111111001111010;
      13'b1110011011100:
        _o_sv = 15'b111111001111011;
      13'b1110011011101:
        _o_sv = 15'b111111001111100;
      13'b1110011011110:
        _o_sv = 15'b111111001111101;
      13'b1110011011111:
        _o_sv = 15'b111111001111110;
      13'b1110011100000:
        _o_sv = 15'b111111001111111;
      13'b1110011100001:
        _o_sv = 15'b111111010000000;
      13'b1110011100010:
        _o_sv = 15'b111111010000001;
      13'b1110011100011:
        _o_sv = 15'b111111010000010;
      13'b1110011100100:
        _o_sv = 15'b111111010000011;
      13'b1110011100101:
        _o_sv = 15'b111111010000100;
      13'b1110011100110:
        _o_sv = 15'b111111010000100;
      13'b1110011100111:
        _o_sv = 15'b111111010000101;
      13'b1110011101000:
        _o_sv = 15'b111111010000110;
      13'b1110011101001:
        _o_sv = 15'b111111010000111;
      13'b1110011101010:
        _o_sv = 15'b111111010001000;
      13'b1110011101011:
        _o_sv = 15'b111111010001001;
      13'b1110011101100:
        _o_sv = 15'b111111010001010;
      13'b1110011101101:
        _o_sv = 15'b111111010001011;
      13'b1110011101110:
        _o_sv = 15'b111111010001100;
      13'b1110011101111:
        _o_sv = 15'b111111010001101;
      13'b1110011110000:
        _o_sv = 15'b111111010001110;
      13'b1110011110001:
        _o_sv = 15'b111111010001111;
      13'b1110011110010:
        _o_sv = 15'b111111010010000;
      13'b1110011110011:
        _o_sv = 15'b111111010010001;
      13'b1110011110100:
        _o_sv = 15'b111111010010010;
      13'b1110011110101:
        _o_sv = 15'b111111010010011;
      13'b1110011110110:
        _o_sv = 15'b111111010010100;
      13'b1110011110111:
        _o_sv = 15'b111111010010100;
      13'b1110011111000:
        _o_sv = 15'b111111010010101;
      13'b1110011111001:
        _o_sv = 15'b111111010010110;
      13'b1110011111010:
        _o_sv = 15'b111111010010111;
      13'b1110011111011:
        _o_sv = 15'b111111010011000;
      13'b1110011111100:
        _o_sv = 15'b111111010011001;
      13'b1110011111101:
        _o_sv = 15'b111111010011010;
      13'b1110011111110:
        _o_sv = 15'b111111010011011;
      13'b1110011111111:
        _o_sv = 15'b111111010011100;
      13'b1110100000000:
        _o_sv = 15'b111111010011101;
      13'b1110100000001:
        _o_sv = 15'b111111010011110;
      13'b1110100000010:
        _o_sv = 15'b111111010011111;
      13'b1110100000011:
        _o_sv = 15'b111111010100000;
      13'b1110100000100:
        _o_sv = 15'b111111010100001;
      13'b1110100000101:
        _o_sv = 15'b111111010100001;
      13'b1110100000110:
        _o_sv = 15'b111111010100010;
      13'b1110100000111:
        _o_sv = 15'b111111010100011;
      13'b1110100001000:
        _o_sv = 15'b111111010100100;
      13'b1110100001001:
        _o_sv = 15'b111111010100101;
      13'b1110100001010:
        _o_sv = 15'b111111010100110;
      13'b1110100001011:
        _o_sv = 15'b111111010100111;
      13'b1110100001100:
        _o_sv = 15'b111111010101000;
      13'b1110100001101:
        _o_sv = 15'b111111010101001;
      13'b1110100001110:
        _o_sv = 15'b111111010101010;
      13'b1110100001111:
        _o_sv = 15'b111111010101011;
      13'b1110100010000:
        _o_sv = 15'b111111010101011;
      13'b1110100010001:
        _o_sv = 15'b111111010101100;
      13'b1110100010010:
        _o_sv = 15'b111111010101101;
      13'b1110100010011:
        _o_sv = 15'b111111010101110;
      13'b1110100010100:
        _o_sv = 15'b111111010101111;
      13'b1110100010101:
        _o_sv = 15'b111111010110000;
      13'b1110100010110:
        _o_sv = 15'b111111010110001;
      13'b1110100010111:
        _o_sv = 15'b111111010110010;
      13'b1110100011000:
        _o_sv = 15'b111111010110011;
      13'b1110100011001:
        _o_sv = 15'b111111010110100;
      13'b1110100011010:
        _o_sv = 15'b111111010110100;
      13'b1110100011011:
        _o_sv = 15'b111111010110101;
      13'b1110100011100:
        _o_sv = 15'b111111010110110;
      13'b1110100011101:
        _o_sv = 15'b111111010110111;
      13'b1110100011110:
        _o_sv = 15'b111111010111000;
      13'b1110100011111:
        _o_sv = 15'b111111010111001;
      13'b1110100100000:
        _o_sv = 15'b111111010111010;
      13'b1110100100001:
        _o_sv = 15'b111111010111011;
      13'b1110100100010:
        _o_sv = 15'b111111010111011;
      13'b1110100100011:
        _o_sv = 15'b111111010111100;
      13'b1110100100100:
        _o_sv = 15'b111111010111101;
      13'b1110100100101:
        _o_sv = 15'b111111010111110;
      13'b1110100100110:
        _o_sv = 15'b111111010111111;
      13'b1110100100111:
        _o_sv = 15'b111111011000000;
      13'b1110100101000:
        _o_sv = 15'b111111011000001;
      13'b1110100101001:
        _o_sv = 15'b111111011000010;
      13'b1110100101010:
        _o_sv = 15'b111111011000011;
      13'b1110100101011:
        _o_sv = 15'b111111011000011;
      13'b1110100101100:
        _o_sv = 15'b111111011000100;
      13'b1110100101101:
        _o_sv = 15'b111111011000101;
      13'b1110100101110:
        _o_sv = 15'b111111011000110;
      13'b1110100101111:
        _o_sv = 15'b111111011000111;
      13'b1110100110000:
        _o_sv = 15'b111111011001000;
      13'b1110100110001:
        _o_sv = 15'b111111011001001;
      13'b1110100110010:
        _o_sv = 15'b111111011001001;
      13'b1110100110011:
        _o_sv = 15'b111111011001010;
      13'b1110100110100:
        _o_sv = 15'b111111011001011;
      13'b1110100110101:
        _o_sv = 15'b111111011001100;
      13'b1110100110110:
        _o_sv = 15'b111111011001101;
      13'b1110100110111:
        _o_sv = 15'b111111011001110;
      13'b1110100111000:
        _o_sv = 15'b111111011001111;
      13'b1110100111001:
        _o_sv = 15'b111111011001111;
      13'b1110100111010:
        _o_sv = 15'b111111011010000;
      13'b1110100111011:
        _o_sv = 15'b111111011010001;
      13'b1110100111100:
        _o_sv = 15'b111111011010010;
      13'b1110100111101:
        _o_sv = 15'b111111011010011;
      13'b1110100111110:
        _o_sv = 15'b111111011010100;
      13'b1110100111111:
        _o_sv = 15'b111111011010101;
      13'b1110101000000:
        _o_sv = 15'b111111011010101;
      13'b1110101000001:
        _o_sv = 15'b111111011010110;
      13'b1110101000010:
        _o_sv = 15'b111111011010111;
      13'b1110101000011:
        _o_sv = 15'b111111011011000;
      13'b1110101000100:
        _o_sv = 15'b111111011011001;
      13'b1110101000101:
        _o_sv = 15'b111111011011010;
      13'b1110101000110:
        _o_sv = 15'b111111011011010;
      13'b1110101000111:
        _o_sv = 15'b111111011011011;
      13'b1110101001000:
        _o_sv = 15'b111111011011100;
      13'b1110101001001:
        _o_sv = 15'b111111011011101;
      13'b1110101001010:
        _o_sv = 15'b111111011011110;
      13'b1110101001011:
        _o_sv = 15'b111111011011111;
      13'b1110101001100:
        _o_sv = 15'b111111011011111;
      13'b1110101001101:
        _o_sv = 15'b111111011100000;
      13'b1110101001110:
        _o_sv = 15'b111111011100001;
      13'b1110101001111:
        _o_sv = 15'b111111011100010;
      13'b1110101010000:
        _o_sv = 15'b111111011100011;
      13'b1110101010001:
        _o_sv = 15'b111111011100100;
      13'b1110101010010:
        _o_sv = 15'b111111011100100;
      13'b1110101010011:
        _o_sv = 15'b111111011100101;
      13'b1110101010100:
        _o_sv = 15'b111111011100110;
      13'b1110101010101:
        _o_sv = 15'b111111011100111;
      13'b1110101010110:
        _o_sv = 15'b111111011101000;
      13'b1110101010111:
        _o_sv = 15'b111111011101001;
      13'b1110101011000:
        _o_sv = 15'b111111011101001;
      13'b1110101011001:
        _o_sv = 15'b111111011101010;
      13'b1110101011010:
        _o_sv = 15'b111111011101011;
      13'b1110101011011:
        _o_sv = 15'b111111011101100;
      13'b1110101011100:
        _o_sv = 15'b111111011101101;
      13'b1110101011101:
        _o_sv = 15'b111111011101101;
      13'b1110101011110:
        _o_sv = 15'b111111011101110;
      13'b1110101011111:
        _o_sv = 15'b111111011101111;
      13'b1110101100000:
        _o_sv = 15'b111111011110000;
      13'b1110101100001:
        _o_sv = 15'b111111011110001;
      13'b1110101100010:
        _o_sv = 15'b111111011110001;
      13'b1110101100011:
        _o_sv = 15'b111111011110010;
      13'b1110101100100:
        _o_sv = 15'b111111011110011;
      13'b1110101100101:
        _o_sv = 15'b111111011110100;
      13'b1110101100110:
        _o_sv = 15'b111111011110101;
      13'b1110101100111:
        _o_sv = 15'b111111011110101;
      13'b1110101101000:
        _o_sv = 15'b111111011110110;
      13'b1110101101001:
        _o_sv = 15'b111111011110111;
      13'b1110101101010:
        _o_sv = 15'b111111011111000;
      13'b1110101101011:
        _o_sv = 15'b111111011111001;
      13'b1110101101100:
        _o_sv = 15'b111111011111001;
      13'b1110101101101:
        _o_sv = 15'b111111011111010;
      13'b1110101101110:
        _o_sv = 15'b111111011111011;
      13'b1110101101111:
        _o_sv = 15'b111111011111100;
      13'b1110101110000:
        _o_sv = 15'b111111011111101;
      13'b1110101110001:
        _o_sv = 15'b111111011111101;
      13'b1110101110010:
        _o_sv = 15'b111111011111110;
      13'b1110101110011:
        _o_sv = 15'b111111011111111;
      13'b1110101110100:
        _o_sv = 15'b111111100000000;
      13'b1110101110101:
        _o_sv = 15'b111111100000001;
      13'b1110101110110:
        _o_sv = 15'b111111100000001;
      13'b1110101110111:
        _o_sv = 15'b111111100000010;
      13'b1110101111000:
        _o_sv = 15'b111111100000011;
      13'b1110101111001:
        _o_sv = 15'b111111100000100;
      13'b1110101111010:
        _o_sv = 15'b111111100000100;
      13'b1110101111011:
        _o_sv = 15'b111111100000101;
      13'b1110101111100:
        _o_sv = 15'b111111100000110;
      13'b1110101111101:
        _o_sv = 15'b111111100000111;
      13'b1110101111110:
        _o_sv = 15'b111111100001000;
      13'b1110101111111:
        _o_sv = 15'b111111100001000;
      13'b1110110000000:
        _o_sv = 15'b111111100001001;
      13'b1110110000001:
        _o_sv = 15'b111111100001010;
      13'b1110110000010:
        _o_sv = 15'b111111100001011;
      13'b1110110000011:
        _o_sv = 15'b111111100001011;
      13'b1110110000100:
        _o_sv = 15'b111111100001100;
      13'b1110110000101:
        _o_sv = 15'b111111100001101;
      13'b1110110000110:
        _o_sv = 15'b111111100001110;
      13'b1110110000111:
        _o_sv = 15'b111111100001110;
      13'b1110110001000:
        _o_sv = 15'b111111100001111;
      13'b1110110001001:
        _o_sv = 15'b111111100010000;
      13'b1110110001010:
        _o_sv = 15'b111111100010001;
      13'b1110110001011:
        _o_sv = 15'b111111100010001;
      13'b1110110001100:
        _o_sv = 15'b111111100010010;
      13'b1110110001101:
        _o_sv = 15'b111111100010011;
      13'b1110110001110:
        _o_sv = 15'b111111100010100;
      13'b1110110001111:
        _o_sv = 15'b111111100010100;
      13'b1110110010000:
        _o_sv = 15'b111111100010101;
      13'b1110110010001:
        _o_sv = 15'b111111100010110;
      13'b1110110010010:
        _o_sv = 15'b111111100010111;
      13'b1110110010011:
        _o_sv = 15'b111111100010111;
      13'b1110110010100:
        _o_sv = 15'b111111100011000;
      13'b1110110010101:
        _o_sv = 15'b111111100011001;
      13'b1110110010110:
        _o_sv = 15'b111111100011010;
      13'b1110110010111:
        _o_sv = 15'b111111100011010;
      13'b1110110011000:
        _o_sv = 15'b111111100011011;
      13'b1110110011001:
        _o_sv = 15'b111111100011100;
      13'b1110110011010:
        _o_sv = 15'b111111100011101;
      13'b1110110011011:
        _o_sv = 15'b111111100011101;
      13'b1110110011100:
        _o_sv = 15'b111111100011110;
      13'b1110110011101:
        _o_sv = 15'b111111100011111;
      13'b1110110011110:
        _o_sv = 15'b111111100100000;
      13'b1110110011111:
        _o_sv = 15'b111111100100000;
      13'b1110110100000:
        _o_sv = 15'b111111100100001;
      13'b1110110100001:
        _o_sv = 15'b111111100100010;
      13'b1110110100010:
        _o_sv = 15'b111111100100011;
      13'b1110110100011:
        _o_sv = 15'b111111100100011;
      13'b1110110100100:
        _o_sv = 15'b111111100100100;
      13'b1110110100101:
        _o_sv = 15'b111111100100101;
      13'b1110110100110:
        _o_sv = 15'b111111100100101;
      13'b1110110100111:
        _o_sv = 15'b111111100100110;
      13'b1110110101000:
        _o_sv = 15'b111111100100111;
      13'b1110110101001:
        _o_sv = 15'b111111100101000;
      13'b1110110101010:
        _o_sv = 15'b111111100101000;
      13'b1110110101011:
        _o_sv = 15'b111111100101001;
      13'b1110110101100:
        _o_sv = 15'b111111100101010;
      13'b1110110101101:
        _o_sv = 15'b111111100101010;
      13'b1110110101110:
        _o_sv = 15'b111111100101011;
      13'b1110110101111:
        _o_sv = 15'b111111100101100;
      13'b1110110110000:
        _o_sv = 15'b111111100101101;
      13'b1110110110001:
        _o_sv = 15'b111111100101101;
      13'b1110110110010:
        _o_sv = 15'b111111100101110;
      13'b1110110110011:
        _o_sv = 15'b111111100101111;
      13'b1110110110100:
        _o_sv = 15'b111111100101111;
      13'b1110110110101:
        _o_sv = 15'b111111100110000;
      13'b1110110110110:
        _o_sv = 15'b111111100110001;
      13'b1110110110111:
        _o_sv = 15'b111111100110010;
      13'b1110110111000:
        _o_sv = 15'b111111100110010;
      13'b1110110111001:
        _o_sv = 15'b111111100110011;
      13'b1110110111010:
        _o_sv = 15'b111111100110100;
      13'b1110110111011:
        _o_sv = 15'b111111100110100;
      13'b1110110111100:
        _o_sv = 15'b111111100110101;
      13'b1110110111101:
        _o_sv = 15'b111111100110110;
      13'b1110110111110:
        _o_sv = 15'b111111100110110;
      13'b1110110111111:
        _o_sv = 15'b111111100110111;
      13'b1110111000000:
        _o_sv = 15'b111111100111000;
      13'b1110111000001:
        _o_sv = 15'b111111100111001;
      13'b1110111000010:
        _o_sv = 15'b111111100111001;
      13'b1110111000011:
        _o_sv = 15'b111111100111010;
      13'b1110111000100:
        _o_sv = 15'b111111100111011;
      13'b1110111000101:
        _o_sv = 15'b111111100111011;
      13'b1110111000110:
        _o_sv = 15'b111111100111100;
      13'b1110111000111:
        _o_sv = 15'b111111100111101;
      13'b1110111001000:
        _o_sv = 15'b111111100111101;
      13'b1110111001001:
        _o_sv = 15'b111111100111110;
      13'b1110111001010:
        _o_sv = 15'b111111100111111;
      13'b1110111001011:
        _o_sv = 15'b111111100111111;
      13'b1110111001100:
        _o_sv = 15'b111111101000000;
      13'b1110111001101:
        _o_sv = 15'b111111101000001;
      13'b1110111001110:
        _o_sv = 15'b111111101000001;
      13'b1110111001111:
        _o_sv = 15'b111111101000010;
      13'b1110111010000:
        _o_sv = 15'b111111101000011;
      13'b1110111010001:
        _o_sv = 15'b111111101000011;
      13'b1110111010010:
        _o_sv = 15'b111111101000100;
      13'b1110111010011:
        _o_sv = 15'b111111101000101;
      13'b1110111010100:
        _o_sv = 15'b111111101000101;
      13'b1110111010101:
        _o_sv = 15'b111111101000110;
      13'b1110111010110:
        _o_sv = 15'b111111101000111;
      13'b1110111010111:
        _o_sv = 15'b111111101000111;
      13'b1110111011000:
        _o_sv = 15'b111111101001000;
      13'b1110111011001:
        _o_sv = 15'b111111101001001;
      13'b1110111011010:
        _o_sv = 15'b111111101001001;
      13'b1110111011011:
        _o_sv = 15'b111111101001010;
      13'b1110111011100:
        _o_sv = 15'b111111101001011;
      13'b1110111011101:
        _o_sv = 15'b111111101001011;
      13'b1110111011110:
        _o_sv = 15'b111111101001100;
      13'b1110111011111:
        _o_sv = 15'b111111101001101;
      13'b1110111100000:
        _o_sv = 15'b111111101001101;
      13'b1110111100001:
        _o_sv = 15'b111111101001110;
      13'b1110111100010:
        _o_sv = 15'b111111101001111;
      13'b1110111100011:
        _o_sv = 15'b111111101001111;
      13'b1110111100100:
        _o_sv = 15'b111111101010000;
      13'b1110111100101:
        _o_sv = 15'b111111101010001;
      13'b1110111100110:
        _o_sv = 15'b111111101010001;
      13'b1110111100111:
        _o_sv = 15'b111111101010010;
      13'b1110111101000:
        _o_sv = 15'b111111101010011;
      13'b1110111101001:
        _o_sv = 15'b111111101010011;
      13'b1110111101010:
        _o_sv = 15'b111111101010100;
      13'b1110111101011:
        _o_sv = 15'b111111101010101;
      13'b1110111101100:
        _o_sv = 15'b111111101010101;
      13'b1110111101101:
        _o_sv = 15'b111111101010110;
      13'b1110111101110:
        _o_sv = 15'b111111101010110;
      13'b1110111101111:
        _o_sv = 15'b111111101010111;
      13'b1110111110000:
        _o_sv = 15'b111111101011000;
      13'b1110111110001:
        _o_sv = 15'b111111101011000;
      13'b1110111110010:
        _o_sv = 15'b111111101011001;
      13'b1110111110011:
        _o_sv = 15'b111111101011010;
      13'b1110111110100:
        _o_sv = 15'b111111101011010;
      13'b1110111110101:
        _o_sv = 15'b111111101011011;
      13'b1110111110110:
        _o_sv = 15'b111111101011011;
      13'b1110111110111:
        _o_sv = 15'b111111101011100;
      13'b1110111111000:
        _o_sv = 15'b111111101011101;
      13'b1110111111001:
        _o_sv = 15'b111111101011101;
      13'b1110111111010:
        _o_sv = 15'b111111101011110;
      13'b1110111111011:
        _o_sv = 15'b111111101011111;
      13'b1110111111100:
        _o_sv = 15'b111111101011111;
      13'b1110111111101:
        _o_sv = 15'b111111101100000;
      13'b1110111111110:
        _o_sv = 15'b111111101100000;
      13'b1110111111111:
        _o_sv = 15'b111111101100001;
      13'b1111000000000:
        _o_sv = 15'b111111101100010;
      13'b1111000000001:
        _o_sv = 15'b111111101100010;
      13'b1111000000010:
        _o_sv = 15'b111111101100011;
      13'b1111000000011:
        _o_sv = 15'b111111101100100;
      13'b1111000000100:
        _o_sv = 15'b111111101100100;
      13'b1111000000101:
        _o_sv = 15'b111111101100101;
      13'b1111000000110:
        _o_sv = 15'b111111101100101;
      13'b1111000000111:
        _o_sv = 15'b111111101100110;
      13'b1111000001000:
        _o_sv = 15'b111111101100111;
      13'b1111000001001:
        _o_sv = 15'b111111101100111;
      13'b1111000001010:
        _o_sv = 15'b111111101101000;
      13'b1111000001011:
        _o_sv = 15'b111111101101000;
      13'b1111000001100:
        _o_sv = 15'b111111101101001;
      13'b1111000001101:
        _o_sv = 15'b111111101101010;
      13'b1111000001110:
        _o_sv = 15'b111111101101010;
      13'b1111000001111:
        _o_sv = 15'b111111101101011;
      13'b1111000010000:
        _o_sv = 15'b111111101101011;
      13'b1111000010001:
        _o_sv = 15'b111111101101100;
      13'b1111000010010:
        _o_sv = 15'b111111101101101;
      13'b1111000010011:
        _o_sv = 15'b111111101101101;
      13'b1111000010100:
        _o_sv = 15'b111111101101110;
      13'b1111000010101:
        _o_sv = 15'b111111101101110;
      13'b1111000010110:
        _o_sv = 15'b111111101101111;
      13'b1111000010111:
        _o_sv = 15'b111111101110000;
      13'b1111000011000:
        _o_sv = 15'b111111101110000;
      13'b1111000011001:
        _o_sv = 15'b111111101110001;
      13'b1111000011010:
        _o_sv = 15'b111111101110001;
      13'b1111000011011:
        _o_sv = 15'b111111101110010;
      13'b1111000011100:
        _o_sv = 15'b111111101110010;
      13'b1111000011101:
        _o_sv = 15'b111111101110011;
      13'b1111000011110:
        _o_sv = 15'b111111101110100;
      13'b1111000011111:
        _o_sv = 15'b111111101110100;
      13'b1111000100000:
        _o_sv = 15'b111111101110101;
      13'b1111000100001:
        _o_sv = 15'b111111101110101;
      13'b1111000100010:
        _o_sv = 15'b111111101110110;
      13'b1111000100011:
        _o_sv = 15'b111111101110111;
      13'b1111000100100:
        _o_sv = 15'b111111101110111;
      13'b1111000100101:
        _o_sv = 15'b111111101111000;
      13'b1111000100110:
        _o_sv = 15'b111111101111000;
      13'b1111000100111:
        _o_sv = 15'b111111101111001;
      13'b1111000101000:
        _o_sv = 15'b111111101111001;
      13'b1111000101001:
        _o_sv = 15'b111111101111010;
      13'b1111000101010:
        _o_sv = 15'b111111101111011;
      13'b1111000101011:
        _o_sv = 15'b111111101111011;
      13'b1111000101100:
        _o_sv = 15'b111111101111100;
      13'b1111000101101:
        _o_sv = 15'b111111101111100;
      13'b1111000101110:
        _o_sv = 15'b111111101111101;
      13'b1111000101111:
        _o_sv = 15'b111111101111101;
      13'b1111000110000:
        _o_sv = 15'b111111101111110;
      13'b1111000110001:
        _o_sv = 15'b111111101111110;
      13'b1111000110010:
        _o_sv = 15'b111111101111111;
      13'b1111000110011:
        _o_sv = 15'b111111110000000;
      13'b1111000110100:
        _o_sv = 15'b111111110000000;
      13'b1111000110101:
        _o_sv = 15'b111111110000001;
      13'b1111000110110:
        _o_sv = 15'b111111110000001;
      13'b1111000110111:
        _o_sv = 15'b111111110000010;
      13'b1111000111000:
        _o_sv = 15'b111111110000010;
      13'b1111000111001:
        _o_sv = 15'b111111110000011;
      13'b1111000111010:
        _o_sv = 15'b111111110000011;
      13'b1111000111011:
        _o_sv = 15'b111111110000100;
      13'b1111000111100:
        _o_sv = 15'b111111110000101;
      13'b1111000111101:
        _o_sv = 15'b111111110000101;
      13'b1111000111110:
        _o_sv = 15'b111111110000110;
      13'b1111000111111:
        _o_sv = 15'b111111110000110;
      13'b1111001000000:
        _o_sv = 15'b111111110000111;
      13'b1111001000001:
        _o_sv = 15'b111111110000111;
      13'b1111001000010:
        _o_sv = 15'b111111110001000;
      13'b1111001000011:
        _o_sv = 15'b111111110001000;
      13'b1111001000100:
        _o_sv = 15'b111111110001001;
      13'b1111001000101:
        _o_sv = 15'b111111110001001;
      13'b1111001000110:
        _o_sv = 15'b111111110001010;
      13'b1111001000111:
        _o_sv = 15'b111111110001010;
      13'b1111001001000:
        _o_sv = 15'b111111110001011;
      13'b1111001001001:
        _o_sv = 15'b111111110001011;
      13'b1111001001010:
        _o_sv = 15'b111111110001100;
      13'b1111001001011:
        _o_sv = 15'b111111110001101;
      13'b1111001001100:
        _o_sv = 15'b111111110001101;
      13'b1111001001101:
        _o_sv = 15'b111111110001110;
      13'b1111001001110:
        _o_sv = 15'b111111110001110;
      13'b1111001001111:
        _o_sv = 15'b111111110001111;
      13'b1111001010000:
        _o_sv = 15'b111111110001111;
      13'b1111001010001:
        _o_sv = 15'b111111110010000;
      13'b1111001010010:
        _o_sv = 15'b111111110010000;
      13'b1111001010011:
        _o_sv = 15'b111111110010001;
      13'b1111001010100:
        _o_sv = 15'b111111110010001;
      13'b1111001010101:
        _o_sv = 15'b111111110010010;
      13'b1111001010110:
        _o_sv = 15'b111111110010010;
      13'b1111001010111:
        _o_sv = 15'b111111110010011;
      13'b1111001011000:
        _o_sv = 15'b111111110010011;
      13'b1111001011001:
        _o_sv = 15'b111111110010100;
      13'b1111001011010:
        _o_sv = 15'b111111110010100;
      13'b1111001011011:
        _o_sv = 15'b111111110010101;
      13'b1111001011100:
        _o_sv = 15'b111111110010101;
      13'b1111001011101:
        _o_sv = 15'b111111110010110;
      13'b1111001011110:
        _o_sv = 15'b111111110010110;
      13'b1111001011111:
        _o_sv = 15'b111111110010111;
      13'b1111001100000:
        _o_sv = 15'b111111110010111;
      13'b1111001100001:
        _o_sv = 15'b111111110011000;
      13'b1111001100010:
        _o_sv = 15'b111111110011000;
      13'b1111001100011:
        _o_sv = 15'b111111110011001;
      13'b1111001100100:
        _o_sv = 15'b111111110011001;
      13'b1111001100101:
        _o_sv = 15'b111111110011010;
      13'b1111001100110:
        _o_sv = 15'b111111110011010;
      13'b1111001100111:
        _o_sv = 15'b111111110011011;
      13'b1111001101000:
        _o_sv = 15'b111111110011011;
      13'b1111001101001:
        _o_sv = 15'b111111110011100;
      13'b1111001101010:
        _o_sv = 15'b111111110011100;
      13'b1111001101011:
        _o_sv = 15'b111111110011101;
      13'b1111001101100:
        _o_sv = 15'b111111110011101;
      13'b1111001101101:
        _o_sv = 15'b111111110011110;
      13'b1111001101110:
        _o_sv = 15'b111111110011110;
      13'b1111001101111:
        _o_sv = 15'b111111110011111;
      13'b1111001110000:
        _o_sv = 15'b111111110011111;
      13'b1111001110001:
        _o_sv = 15'b111111110100000;
      13'b1111001110010:
        _o_sv = 15'b111111110100000;
      13'b1111001110011:
        _o_sv = 15'b111111110100001;
      13'b1111001110100:
        _o_sv = 15'b111111110100001;
      13'b1111001110101:
        _o_sv = 15'b111111110100010;
      13'b1111001110110:
        _o_sv = 15'b111111110100010;
      13'b1111001110111:
        _o_sv = 15'b111111110100011;
      13'b1111001111000:
        _o_sv = 15'b111111110100011;
      13'b1111001111001:
        _o_sv = 15'b111111110100011;
      13'b1111001111010:
        _o_sv = 15'b111111110100100;
      13'b1111001111011:
        _o_sv = 15'b111111110100100;
      13'b1111001111100:
        _o_sv = 15'b111111110100101;
      13'b1111001111101:
        _o_sv = 15'b111111110100101;
      13'b1111001111110:
        _o_sv = 15'b111111110100110;
      13'b1111001111111:
        _o_sv = 15'b111111110100110;
      13'b1111010000000:
        _o_sv = 15'b111111110100111;
      13'b1111010000001:
        _o_sv = 15'b111111110100111;
      13'b1111010000010:
        _o_sv = 15'b111111110101000;
      13'b1111010000011:
        _o_sv = 15'b111111110101000;
      13'b1111010000100:
        _o_sv = 15'b111111110101001;
      13'b1111010000101:
        _o_sv = 15'b111111110101001;
      13'b1111010000110:
        _o_sv = 15'b111111110101001;
      13'b1111010000111:
        _o_sv = 15'b111111110101010;
      13'b1111010001000:
        _o_sv = 15'b111111110101010;
      13'b1111010001001:
        _o_sv = 15'b111111110101011;
      13'b1111010001010:
        _o_sv = 15'b111111110101011;
      13'b1111010001011:
        _o_sv = 15'b111111110101100;
      13'b1111010001100:
        _o_sv = 15'b111111110101100;
      13'b1111010001101:
        _o_sv = 15'b111111110101101;
      13'b1111010001110:
        _o_sv = 15'b111111110101101;
      13'b1111010001111:
        _o_sv = 15'b111111110101110;
      13'b1111010010000:
        _o_sv = 15'b111111110101110;
      13'b1111010010001:
        _o_sv = 15'b111111110101110;
      13'b1111010010010:
        _o_sv = 15'b111111110101111;
      13'b1111010010011:
        _o_sv = 15'b111111110101111;
      13'b1111010010100:
        _o_sv = 15'b111111110110000;
      13'b1111010010101:
        _o_sv = 15'b111111110110000;
      13'b1111010010110:
        _o_sv = 15'b111111110110001;
      13'b1111010010111:
        _o_sv = 15'b111111110110001;
      13'b1111010011000:
        _o_sv = 15'b111111110110001;
      13'b1111010011001:
        _o_sv = 15'b111111110110010;
      13'b1111010011010:
        _o_sv = 15'b111111110110010;
      13'b1111010011011:
        _o_sv = 15'b111111110110011;
      13'b1111010011100:
        _o_sv = 15'b111111110110011;
      13'b1111010011101:
        _o_sv = 15'b111111110110100;
      13'b1111010011110:
        _o_sv = 15'b111111110110100;
      13'b1111010011111:
        _o_sv = 15'b111111110110100;
      13'b1111010100000:
        _o_sv = 15'b111111110110101;
      13'b1111010100001:
        _o_sv = 15'b111111110110101;
      13'b1111010100010:
        _o_sv = 15'b111111110110110;
      13'b1111010100011:
        _o_sv = 15'b111111110110110;
      13'b1111010100100:
        _o_sv = 15'b111111110110111;
      13'b1111010100101:
        _o_sv = 15'b111111110110111;
      13'b1111010100110:
        _o_sv = 15'b111111110110111;
      13'b1111010100111:
        _o_sv = 15'b111111110111000;
      13'b1111010101000:
        _o_sv = 15'b111111110111000;
      13'b1111010101001:
        _o_sv = 15'b111111110111001;
      13'b1111010101010:
        _o_sv = 15'b111111110111001;
      13'b1111010101011:
        _o_sv = 15'b111111110111001;
      13'b1111010101100:
        _o_sv = 15'b111111110111010;
      13'b1111010101101:
        _o_sv = 15'b111111110111010;
      13'b1111010101110:
        _o_sv = 15'b111111110111011;
      13'b1111010101111:
        _o_sv = 15'b111111110111011;
      13'b1111010110000:
        _o_sv = 15'b111111110111100;
      13'b1111010110001:
        _o_sv = 15'b111111110111100;
      13'b1111010110010:
        _o_sv = 15'b111111110111100;
      13'b1111010110011:
        _o_sv = 15'b111111110111101;
      13'b1111010110100:
        _o_sv = 15'b111111110111101;
      13'b1111010110101:
        _o_sv = 15'b111111110111110;
      13'b1111010110110:
        _o_sv = 15'b111111110111110;
      13'b1111010110111:
        _o_sv = 15'b111111110111110;
      13'b1111010111000:
        _o_sv = 15'b111111110111111;
      13'b1111010111001:
        _o_sv = 15'b111111110111111;
      13'b1111010111010:
        _o_sv = 15'b111111111000000;
      13'b1111010111011:
        _o_sv = 15'b111111111000000;
      13'b1111010111100:
        _o_sv = 15'b111111111000000;
      13'b1111010111101:
        _o_sv = 15'b111111111000001;
      13'b1111010111110:
        _o_sv = 15'b111111111000001;
      13'b1111010111111:
        _o_sv = 15'b111111111000001;
      13'b1111011000000:
        _o_sv = 15'b111111111000010;
      13'b1111011000001:
        _o_sv = 15'b111111111000010;
      13'b1111011000010:
        _o_sv = 15'b111111111000011;
      13'b1111011000011:
        _o_sv = 15'b111111111000011;
      13'b1111011000100:
        _o_sv = 15'b111111111000011;
      13'b1111011000101:
        _o_sv = 15'b111111111000100;
      13'b1111011000110:
        _o_sv = 15'b111111111000100;
      13'b1111011000111:
        _o_sv = 15'b111111111000101;
      13'b1111011001000:
        _o_sv = 15'b111111111000101;
      13'b1111011001001:
        _o_sv = 15'b111111111000101;
      13'b1111011001010:
        _o_sv = 15'b111111111000110;
      13'b1111011001011:
        _o_sv = 15'b111111111000110;
      13'b1111011001100:
        _o_sv = 15'b111111111000110;
      13'b1111011001101:
        _o_sv = 15'b111111111000111;
      13'b1111011001110:
        _o_sv = 15'b111111111000111;
      13'b1111011001111:
        _o_sv = 15'b111111111000111;
      13'b1111011010000:
        _o_sv = 15'b111111111001000;
      13'b1111011010001:
        _o_sv = 15'b111111111001000;
      13'b1111011010010:
        _o_sv = 15'b111111111001001;
      13'b1111011010011:
        _o_sv = 15'b111111111001001;
      13'b1111011010100:
        _o_sv = 15'b111111111001001;
      13'b1111011010101:
        _o_sv = 15'b111111111001010;
      13'b1111011010110:
        _o_sv = 15'b111111111001010;
      13'b1111011010111:
        _o_sv = 15'b111111111001010;
      13'b1111011011000:
        _o_sv = 15'b111111111001011;
      13'b1111011011001:
        _o_sv = 15'b111111111001011;
      13'b1111011011010:
        _o_sv = 15'b111111111001011;
      13'b1111011011011:
        _o_sv = 15'b111111111001100;
      13'b1111011011100:
        _o_sv = 15'b111111111001100;
      13'b1111011011101:
        _o_sv = 15'b111111111001101;
      13'b1111011011110:
        _o_sv = 15'b111111111001101;
      13'b1111011011111:
        _o_sv = 15'b111111111001101;
      13'b1111011100000:
        _o_sv = 15'b111111111001110;
      13'b1111011100001:
        _o_sv = 15'b111111111001110;
      13'b1111011100010:
        _o_sv = 15'b111111111001110;
      13'b1111011100011:
        _o_sv = 15'b111111111001111;
      13'b1111011100100:
        _o_sv = 15'b111111111001111;
      13'b1111011100101:
        _o_sv = 15'b111111111001111;
      13'b1111011100110:
        _o_sv = 15'b111111111010000;
      13'b1111011100111:
        _o_sv = 15'b111111111010000;
      13'b1111011101000:
        _o_sv = 15'b111111111010000;
      13'b1111011101001:
        _o_sv = 15'b111111111010001;
      13'b1111011101010:
        _o_sv = 15'b111111111010001;
      13'b1111011101011:
        _o_sv = 15'b111111111010001;
      13'b1111011101100:
        _o_sv = 15'b111111111010010;
      13'b1111011101101:
        _o_sv = 15'b111111111010010;
      13'b1111011101110:
        _o_sv = 15'b111111111010010;
      13'b1111011101111:
        _o_sv = 15'b111111111010011;
      13'b1111011110000:
        _o_sv = 15'b111111111010011;
      13'b1111011110001:
        _o_sv = 15'b111111111010011;
      13'b1111011110010:
        _o_sv = 15'b111111111010100;
      13'b1111011110011:
        _o_sv = 15'b111111111010100;
      13'b1111011110100:
        _o_sv = 15'b111111111010100;
      13'b1111011110101:
        _o_sv = 15'b111111111010101;
      13'b1111011110110:
        _o_sv = 15'b111111111010101;
      13'b1111011110111:
        _o_sv = 15'b111111111010101;
      13'b1111011111000:
        _o_sv = 15'b111111111010110;
      13'b1111011111001:
        _o_sv = 15'b111111111010110;
      13'b1111011111010:
        _o_sv = 15'b111111111010110;
      13'b1111011111011:
        _o_sv = 15'b111111111010110;
      13'b1111011111100:
        _o_sv = 15'b111111111010111;
      13'b1111011111101:
        _o_sv = 15'b111111111010111;
      13'b1111011111110:
        _o_sv = 15'b111111111010111;
      13'b1111011111111:
        _o_sv = 15'b111111111011000;
      13'b1111100000000:
        _o_sv = 15'b111111111011000;
      13'b1111100000001:
        _o_sv = 15'b111111111011000;
      13'b1111100000010:
        _o_sv = 15'b111111111011001;
      13'b1111100000011:
        _o_sv = 15'b111111111011001;
      13'b1111100000100:
        _o_sv = 15'b111111111011001;
      13'b1111100000101:
        _o_sv = 15'b111111111011010;
      13'b1111100000110:
        _o_sv = 15'b111111111011010;
      13'b1111100000111:
        _o_sv = 15'b111111111011010;
      13'b1111100001000:
        _o_sv = 15'b111111111011010;
      13'b1111100001001:
        _o_sv = 15'b111111111011011;
      13'b1111100001010:
        _o_sv = 15'b111111111011011;
      13'b1111100001011:
        _o_sv = 15'b111111111011011;
      13'b1111100001100:
        _o_sv = 15'b111111111011100;
      13'b1111100001101:
        _o_sv = 15'b111111111011100;
      13'b1111100001110:
        _o_sv = 15'b111111111011100;
      13'b1111100001111:
        _o_sv = 15'b111111111011101;
      13'b1111100010000:
        _o_sv = 15'b111111111011101;
      13'b1111100010001:
        _o_sv = 15'b111111111011101;
      13'b1111100010010:
        _o_sv = 15'b111111111011101;
      13'b1111100010011:
        _o_sv = 15'b111111111011110;
      13'b1111100010100:
        _o_sv = 15'b111111111011110;
      13'b1111100010101:
        _o_sv = 15'b111111111011110;
      13'b1111100010110:
        _o_sv = 15'b111111111011111;
      13'b1111100010111:
        _o_sv = 15'b111111111011111;
      13'b1111100011000:
        _o_sv = 15'b111111111011111;
      13'b1111100011001:
        _o_sv = 15'b111111111011111;
      13'b1111100011010:
        _o_sv = 15'b111111111100000;
      13'b1111100011011:
        _o_sv = 15'b111111111100000;
      13'b1111100011100:
        _o_sv = 15'b111111111100000;
      13'b1111100011101:
        _o_sv = 15'b111111111100000;
      13'b1111100011110:
        _o_sv = 15'b111111111100001;
      13'b1111100011111:
        _o_sv = 15'b111111111100001;
      13'b1111100100000:
        _o_sv = 15'b111111111100001;
      13'b1111100100001:
        _o_sv = 15'b111111111100010;
      13'b1111100100010:
        _o_sv = 15'b111111111100010;
      13'b1111100100011:
        _o_sv = 15'b111111111100010;
      13'b1111100100100:
        _o_sv = 15'b111111111100010;
      13'b1111100100101:
        _o_sv = 15'b111111111100011;
      13'b1111100100110:
        _o_sv = 15'b111111111100011;
      13'b1111100100111:
        _o_sv = 15'b111111111100011;
      13'b1111100101000:
        _o_sv = 15'b111111111100011;
      13'b1111100101001:
        _o_sv = 15'b111111111100100;
      13'b1111100101010:
        _o_sv = 15'b111111111100100;
      13'b1111100101011:
        _o_sv = 15'b111111111100100;
      13'b1111100101100:
        _o_sv = 15'b111111111100100;
      13'b1111100101101:
        _o_sv = 15'b111111111100101;
      13'b1111100101110:
        _o_sv = 15'b111111111100101;
      13'b1111100101111:
        _o_sv = 15'b111111111100101;
      13'b1111100110000:
        _o_sv = 15'b111111111100101;
      13'b1111100110001:
        _o_sv = 15'b111111111100110;
      13'b1111100110010:
        _o_sv = 15'b111111111100110;
      13'b1111100110011:
        _o_sv = 15'b111111111100110;
      13'b1111100110100:
        _o_sv = 15'b111111111100110;
      13'b1111100110101:
        _o_sv = 15'b111111111100111;
      13'b1111100110110:
        _o_sv = 15'b111111111100111;
      13'b1111100110111:
        _o_sv = 15'b111111111100111;
      13'b1111100111000:
        _o_sv = 15'b111111111100111;
      13'b1111100111001:
        _o_sv = 15'b111111111101000;
      13'b1111100111010:
        _o_sv = 15'b111111111101000;
      13'b1111100111011:
        _o_sv = 15'b111111111101000;
      13'b1111100111100:
        _o_sv = 15'b111111111101000;
      13'b1111100111101:
        _o_sv = 15'b111111111101001;
      13'b1111100111110:
        _o_sv = 15'b111111111101001;
      13'b1111100111111:
        _o_sv = 15'b111111111101001;
      13'b1111101000000:
        _o_sv = 15'b111111111101001;
      13'b1111101000001:
        _o_sv = 15'b111111111101010;
      13'b1111101000010:
        _o_sv = 15'b111111111101010;
      13'b1111101000011:
        _o_sv = 15'b111111111101010;
      13'b1111101000100:
        _o_sv = 15'b111111111101010;
      13'b1111101000101:
        _o_sv = 15'b111111111101010;
      13'b1111101000110:
        _o_sv = 15'b111111111101011;
      13'b1111101000111:
        _o_sv = 15'b111111111101011;
      13'b1111101001000:
        _o_sv = 15'b111111111101011;
      13'b1111101001001:
        _o_sv = 15'b111111111101011;
      13'b1111101001010:
        _o_sv = 15'b111111111101100;
      13'b1111101001011:
        _o_sv = 15'b111111111101100;
      13'b1111101001100:
        _o_sv = 15'b111111111101100;
      13'b1111101001101:
        _o_sv = 15'b111111111101100;
      13'b1111101001110:
        _o_sv = 15'b111111111101100;
      13'b1111101001111:
        _o_sv = 15'b111111111101101;
      13'b1111101010000:
        _o_sv = 15'b111111111101101;
      13'b1111101010001:
        _o_sv = 15'b111111111101101;
      13'b1111101010010:
        _o_sv = 15'b111111111101101;
      13'b1111101010011:
        _o_sv = 15'b111111111101101;
      13'b1111101010100:
        _o_sv = 15'b111111111101110;
      13'b1111101010101:
        _o_sv = 15'b111111111101110;
      13'b1111101010110:
        _o_sv = 15'b111111111101110;
      13'b1111101010111:
        _o_sv = 15'b111111111101110;
      13'b1111101011000:
        _o_sv = 15'b111111111101110;
      13'b1111101011001:
        _o_sv = 15'b111111111101111;
      13'b1111101011010:
        _o_sv = 15'b111111111101111;
      13'b1111101011011:
        _o_sv = 15'b111111111101111;
      13'b1111101011100:
        _o_sv = 15'b111111111101111;
      13'b1111101011101:
        _o_sv = 15'b111111111101111;
      13'b1111101011110:
        _o_sv = 15'b111111111110000;
      13'b1111101011111:
        _o_sv = 15'b111111111110000;
      13'b1111101100000:
        _o_sv = 15'b111111111110000;
      13'b1111101100001:
        _o_sv = 15'b111111111110000;
      13'b1111101100010:
        _o_sv = 15'b111111111110000;
      13'b1111101100011:
        _o_sv = 15'b111111111110001;
      13'b1111101100100:
        _o_sv = 15'b111111111110001;
      13'b1111101100101:
        _o_sv = 15'b111111111110001;
      13'b1111101100110:
        _o_sv = 15'b111111111110001;
      13'b1111101100111:
        _o_sv = 15'b111111111110001;
      13'b1111101101000:
        _o_sv = 15'b111111111110010;
      13'b1111101101001:
        _o_sv = 15'b111111111110010;
      13'b1111101101010:
        _o_sv = 15'b111111111110010;
      13'b1111101101011:
        _o_sv = 15'b111111111110010;
      13'b1111101101100:
        _o_sv = 15'b111111111110010;
      13'b1111101101101:
        _o_sv = 15'b111111111110010;
      13'b1111101101110:
        _o_sv = 15'b111111111110011;
      13'b1111101101111:
        _o_sv = 15'b111111111110011;
      13'b1111101110000:
        _o_sv = 15'b111111111110011;
      13'b1111101110001:
        _o_sv = 15'b111111111110011;
      13'b1111101110010:
        _o_sv = 15'b111111111110011;
      13'b1111101110011:
        _o_sv = 15'b111111111110100;
      13'b1111101110100:
        _o_sv = 15'b111111111110100;
      13'b1111101110101:
        _o_sv = 15'b111111111110100;
      13'b1111101110110:
        _o_sv = 15'b111111111110100;
      13'b1111101110111:
        _o_sv = 15'b111111111110100;
      13'b1111101111000:
        _o_sv = 15'b111111111110100;
      13'b1111101111001:
        _o_sv = 15'b111111111110101;
      13'b1111101111010:
        _o_sv = 15'b111111111110101;
      13'b1111101111011:
        _o_sv = 15'b111111111110101;
      13'b1111101111100:
        _o_sv = 15'b111111111110101;
      13'b1111101111101:
        _o_sv = 15'b111111111110101;
      13'b1111101111110:
        _o_sv = 15'b111111111110101;
      13'b1111101111111:
        _o_sv = 15'b111111111110101;
      13'b1111110000000:
        _o_sv = 15'b111111111110110;
      13'b1111110000001:
        _o_sv = 15'b111111111110110;
      13'b1111110000010:
        _o_sv = 15'b111111111110110;
      13'b1111110000011:
        _o_sv = 15'b111111111110110;
      13'b1111110000100:
        _o_sv = 15'b111111111110110;
      13'b1111110000101:
        _o_sv = 15'b111111111110110;
      13'b1111110000110:
        _o_sv = 15'b111111111110111;
      13'b1111110000111:
        _o_sv = 15'b111111111110111;
      13'b1111110001000:
        _o_sv = 15'b111111111110111;
      13'b1111110001001:
        _o_sv = 15'b111111111110111;
      13'b1111110001010:
        _o_sv = 15'b111111111110111;
      13'b1111110001011:
        _o_sv = 15'b111111111110111;
      13'b1111110001100:
        _o_sv = 15'b111111111110111;
      13'b1111110001101:
        _o_sv = 15'b111111111111000;
      13'b1111110001110:
        _o_sv = 15'b111111111111000;
      13'b1111110001111:
        _o_sv = 15'b111111111111000;
      13'b1111110010000:
        _o_sv = 15'b111111111111000;
      13'b1111110010001:
        _o_sv = 15'b111111111111000;
      13'b1111110010010:
        _o_sv = 15'b111111111111000;
      13'b1111110010011:
        _o_sv = 15'b111111111111000;
      13'b1111110010100:
        _o_sv = 15'b111111111111000;
      13'b1111110010101:
        _o_sv = 15'b111111111111001;
      13'b1111110010110:
        _o_sv = 15'b111111111111001;
      13'b1111110010111:
        _o_sv = 15'b111111111111001;
      13'b1111110011000:
        _o_sv = 15'b111111111111001;
      13'b1111110011001:
        _o_sv = 15'b111111111111001;
      13'b1111110011010:
        _o_sv = 15'b111111111111001;
      13'b1111110011011:
        _o_sv = 15'b111111111111001;
      13'b1111110011100:
        _o_sv = 15'b111111111111001;
      13'b1111110011101:
        _o_sv = 15'b111111111111010;
      13'b1111110011110:
        _o_sv = 15'b111111111111010;
      13'b1111110011111:
        _o_sv = 15'b111111111111010;
      13'b1111110100000:
        _o_sv = 15'b111111111111010;
      13'b1111110100001:
        _o_sv = 15'b111111111111010;
      13'b1111110100010:
        _o_sv = 15'b111111111111010;
      13'b1111110100011:
        _o_sv = 15'b111111111111010;
      13'b1111110100100:
        _o_sv = 15'b111111111111010;
      13'b1111110100101:
        _o_sv = 15'b111111111111011;
      13'b1111110100110:
        _o_sv = 15'b111111111111011;
      13'b1111110100111:
        _o_sv = 15'b111111111111011;
      13'b1111110101000:
        _o_sv = 15'b111111111111011;
      13'b1111110101001:
        _o_sv = 15'b111111111111011;
      13'b1111110101010:
        _o_sv = 15'b111111111111011;
      13'b1111110101011:
        _o_sv = 15'b111111111111011;
      13'b1111110101100:
        _o_sv = 15'b111111111111011;
      13'b1111110101101:
        _o_sv = 15'b111111111111011;
      13'b1111110101110:
        _o_sv = 15'b111111111111011;
      13'b1111110101111:
        _o_sv = 15'b111111111111100;
      13'b1111110110000:
        _o_sv = 15'b111111111111100;
      13'b1111110110001:
        _o_sv = 15'b111111111111100;
      13'b1111110110010:
        _o_sv = 15'b111111111111100;
      13'b1111110110011:
        _o_sv = 15'b111111111111100;
      13'b1111110110100:
        _o_sv = 15'b111111111111100;
      13'b1111110110101:
        _o_sv = 15'b111111111111100;
      13'b1111110110110:
        _o_sv = 15'b111111111111100;
      13'b1111110110111:
        _o_sv = 15'b111111111111100;
      13'b1111110111000:
        _o_sv = 15'b111111111111100;
      13'b1111110111001:
        _o_sv = 15'b111111111111100;
      13'b1111110111010:
        _o_sv = 15'b111111111111101;
      13'b1111110111011:
        _o_sv = 15'b111111111111101;
      13'b1111110111100:
        _o_sv = 15'b111111111111101;
      13'b1111110111101:
        _o_sv = 15'b111111111111101;
      13'b1111110111110:
        _o_sv = 15'b111111111111101;
      13'b1111110111111:
        _o_sv = 15'b111111111111101;
      13'b1111111000000:
        _o_sv = 15'b111111111111101;
      13'b1111111000001:
        _o_sv = 15'b111111111111101;
      13'b1111111000010:
        _o_sv = 15'b111111111111101;
      13'b1111111000011:
        _o_sv = 15'b111111111111101;
      13'b1111111000100:
        _o_sv = 15'b111111111111101;
      13'b1111111000101:
        _o_sv = 15'b111111111111101;
      13'b1111111000110:
        _o_sv = 15'b111111111111101;
      13'b1111111000111:
        _o_sv = 15'b111111111111110;
      13'b1111111001000:
        _o_sv = 15'b111111111111110;
      13'b1111111001001:
        _o_sv = 15'b111111111111110;
      13'b1111111001010:
        _o_sv = 15'b111111111111110;
      13'b1111111001011:
        _o_sv = 15'b111111111111110;
      13'b1111111001100:
        _o_sv = 15'b111111111111110;
      13'b1111111001101:
        _o_sv = 15'b111111111111110;
      13'b1111111001110:
        _o_sv = 15'b111111111111110;
      13'b1111111001111:
        _o_sv = 15'b111111111111110;
      13'b1111111010000:
        _o_sv = 15'b111111111111110;
      13'b1111111010001:
        _o_sv = 15'b111111111111110;
      13'b1111111010010:
        _o_sv = 15'b111111111111110;
      13'b1111111010011:
        _o_sv = 15'b111111111111110;
      13'b1111111010100:
        _o_sv = 15'b111111111111110;
      13'b1111111010101:
        _o_sv = 15'b111111111111110;
      13'b1111111010110:
        _o_sv = 15'b111111111111110;
      13'b1111111010111:
        _o_sv = 15'b111111111111110;
      13'b1111111011000:
        _o_sv = 15'b111111111111111;
      13'b1111111011001:
        _o_sv = 15'b111111111111111;
      13'b1111111011010:
        _o_sv = 15'b111111111111111;
      13'b1111111011011:
        _o_sv = 15'b111111111111111;
      13'b1111111011100:
        _o_sv = 15'b111111111111111;
      13'b1111111011101:
        _o_sv = 15'b111111111111111;
      13'b1111111011110:
        _o_sv = 15'b111111111111111;
      13'b1111111011111:
        _o_sv = 15'b111111111111111;
      13'b1111111100000:
        _o_sv = 15'b111111111111111;
      13'b1111111100001:
        _o_sv = 15'b111111111111111;
      13'b1111111100010:
        _o_sv = 15'b111111111111111;
      13'b1111111100011:
        _o_sv = 15'b111111111111111;
      13'b1111111100100:
        _o_sv = 15'b111111111111111;
      13'b1111111100101:
        _o_sv = 15'b111111111111111;
      13'b1111111100110:
        _o_sv = 15'b111111111111111;
      13'b1111111100111:
        _o_sv = 15'b111111111111111;
      13'b1111111101000:
        _o_sv = 15'b111111111111111;
      13'b1111111101001:
        _o_sv = 15'b111111111111111;
      13'b1111111101010:
        _o_sv = 15'b111111111111111;
      13'b1111111101011:
        _o_sv = 15'b111111111111111;
      13'b1111111101100:
        _o_sv = 15'b111111111111111;
      13'b1111111101101:
        _o_sv = 15'b111111111111111;
      13'b1111111101110:
        _o_sv = 15'b111111111111111;
      13'b1111111101111:
        _o_sv = 15'b111111111111111;
      13'b1111111110000:
        _o_sv = 15'b111111111111111;
      13'b1111111110001:
        _o_sv = 15'b111111111111111;
      13'b1111111110010:
        _o_sv = 15'b111111111111111;
      13'b1111111110011:
        _o_sv = 15'b111111111111111;
      13'b1111111110100:
        _o_sv = 15'b111111111111111;
      13'b1111111110101:
        _o_sv = 15'b111111111111111;
      13'b1111111110110:
        _o_sv = 15'b111111111111111;
      13'b1111111110111:
        _o_sv = 15'b111111111111111;
      13'b1111111111000:
        _o_sv = 15'b111111111111111;
      13'b1111111111001:
        _o_sv = 15'b111111111111111;
      13'b1111111111010:
        _o_sv = 15'b111111111111111;
      13'b1111111111011:
        _o_sv = 15'b111111111111111;
      13'b1111111111100:
        _o_sv = 15'b111111111111111;
      13'b1111111111101:
        _o_sv = 15'b111111111111111;
      13'b1111111111110:
        _o_sv = 15'b111111111111111;
      13'b1111111111111:
        _o_sv = 15'b111111111111111;
    endcase
  end
endmodule // sine
